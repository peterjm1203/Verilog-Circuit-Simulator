
module main(g35,g36,g6744,g6745,g6746,g6747,g6748,g6749,g6750,g6751,g6752,g6753,g84,g120,g5,g113,g126,g99,g53,g116,g92,g56,g91,g44,g57,g100,g54,g124,g125,g114,g134,g72,g115,g135,g90,g127,g64,g73,g7243,g7245,g7257,g7260,g7540,g7916,g7946,g8132,g8178,g8215,g8235,g8277,g8279,g8283,g8291,g8342,g8344,g8353,g8358,g8398,g8403,g8416,g8475,g8719,g8783,g8784,g8785,g8786,g8787,g8788,g8789,g8839,g8870,g8915,g8916,g8917,g8918,g8919,g8920,g9019,g9048,g9251,g9497,g9553,g9555,g9615,g9617,g9680,g9682,g9741,g9743,g9817,g10122,g10306,g10500,g10527,g11349,g11388,g11418,g11447,g11678,g11770,g12184,g12238,g12300,g12350,g12368,g12422,g12470,g12832,g12919,g12923,g13039,g13049,g13068,g13085,g13099,g13259,g13272,g13865,g13881,g13895,g13906,g13926,g13966,g14096,g14125,g14147,g14167,g14189,g14201,g14217,g14421,g14451,g14518,g14597,g14635,g14662,g14673,g14694,g14705,g14738,g14749,g14779,g14828,g16603,g16624,g16627,g16656,g16659,g16686,g16693,g16718,g16722,g16744,g16748,g16775,g16874,g16924,g16955,g17291,g17316,g17320,g17400,g17404,g17423,g17519,g17577,g17580,g17604,g17607,g17639,g17646,g17649,g17674,g17678,g17685,g17688,g17711,g17715,g17722,g17739,g17743,g17760,g17764,g17778,g17787,g17813,g17819,g17845,g17871,g18092,g18094,g18095,g18096,g18097,g18098,g18099,g18100,g18101,g18881,g19334,g19357,g20049,g20557,g20652,g20654,g20763,g20899,g20901,g21176,g21245,g21270,g21292,g21698,g21727,g23002,g23190,g23612,g23652,g23683,g23759,g24151,g25114,g25167,g25219,g25259,g25582,g25583,g25584,g25585,g25586,g25587,g25588,g25589,g25590,g26801,g26875,g26876,g26877,g27831,g28030,g28041,g28042,g28753,g29210,g29211,g29212,g29213,g29214,g29215,g29216,g29217,g29218,g29219,g29220,g29221,g30327,g30329,g30330,g30331,g30332,g31521,g31656,g31665,g31793,g31860,g31861,g31862,g31863,g32185,g32429,g32454,g32975,g33079,g33435,g33533,g33636,g33659,g33874,g33894,g33935,g33945,g33946,g33947,g33948,g33949,g33950,g33959,g34201,g34221,g34232,g34233,g34234,g34235,g34236,g34237,g34238,g34239,g34240,g34383,g34425,g34435,g34436,g34437,g34597,g34788,g34839,g34913,g34915,g34917,g34919,g34921,g34923,g34925,g34927,g34956,g34972,g24168,g24178,g12833,g24174,g24181,g24172,g24161,g24177,g24171,g24163,g24170,g24185,g24164,g24173,g24162,g24179,g24180,g24175,g24183,g24166,g24176,g24184,g24169,g24182,g24165,g24167);

input g35;
input g36;
input g6744;
input g6745;
input g6746;
input g6747;
input g6748;
input g6749;
input g6750;
input g6751;
input g6752;
input g6753;
input g84;
input g120;
input g5;
input g113;
input g126;
input g99;
input g53;
input g116;
input g92;
input g56;
input g91;
input g44;
input g57;
input g100;
input g54;
input g124;
input g125;
input g114;
input g134;
input g72;
input g115;
input g135;
input g90;
input g127;
input g64;
input g73;

output g7243;
output g7245;
output g7257;
output g7260;
output g7540;
output g7916;
output g7946;
output g8132;
output g8178;
output g8215;
output g8235;
output g8277;
output g8279;
output g8283;
output g8291;
output g8342;
output g8344;
output g8353;
output g8358;
output g8398;
output g8403;
output g8416;
output g8475;
output g8719;
output g8783;
output g8784;
output g8785;
output g8786;
output g8787;
output g8788;
output g8789;
output g8839;
output g8870;
output g8915;
output g8916;
output g8917;
output g8918;
output g8919;
output g8920;
output g9019;
output g9048;
output g9251;
output g9497;
output g9553;
output g9555;
output g9615;
output g9617;
output g9680;
output g9682;
output g9741;
output g9743;
output g9817;
output g10122;
output g10306;
output g10500;
output g10527;
output g11349;
output g11388;
output g11418;
output g11447;
output g11678;
output g11770;
output g12184;
output g12238;
output g12300;
output g12350;
output g12368;
output g12422;
output g12470;
output g12832;
output g12919;
output g12923;
output g13039;
output g13049;
output g13068;
output g13085;
output g13099;
output g13259;
output g13272;
output g13865;
output g13881;
output g13895;
output g13906;
output g13926;
output g13966;
output g14096;
output g14125;
output g14147;
output g14167;
output g14189;
output g14201;
output g14217;
output g14421;
output g14451;
output g14518;
output g14597;
output g14635;
output g14662;
output g14673;
output g14694;
output g14705;
output g14738;
output g14749;
output g14779;
output g14828;
output g16603;
output g16624;
output g16627;
output g16656;
output g16659;
output g16686;
output g16693;
output g16718;
output g16722;
output g16744;
output g16748;
output g16775;
output g16874;
output g16924;
output g16955;
output g17291;
output g17316;
output g17320;
output g17400;
output g17404;
output g17423;
output g17519;
output g17577;
output g17580;
output g17604;
output g17607;
output g17639;
output g17646;
output g17649;
output g17674;
output g17678;
output g17685;
output g17688;
output g17711;
output g17715;
output g17722;
output g17739;
output g17743;
output g17760;
output g17764;
output g17778;
output g17787;
output g17813;
output g17819;
output g17845;
output g17871;
output g18092;
output g18094;
output g18095;
output g18096;
output g18097;
output g18098;
output g18099;
output g18100;
output g18101;
output g18881;
output g19334;
output g19357;
output g20049;
output g20557;
output g20652;
output g20654;
output g20763;
output g20899;
output g20901;
output g21176;
output g21245;
output g21270;
output g21292;
output g21698;
output g21727;
output g23002;
output g23190;
output g23612;
output g23652;
output g23683;
output g23759;
output g24151;
output g25114;
output g25167;
output g25219;
output g25259;
output g25582;
output g25583;
output g25584;
output g25585;
output g25586;
output g25587;
output g25588;
output g25589;
output g25590;
output g26801;
output g26875;
output g26876;
output g26877;
output g27831;
output g28030;
output g28041;
output g28042;
output g28753;
output g29210;
output g29211;
output g29212;
output g29213;
output g29214;
output g29215;
output g29216;
output g29217;
output g29218;
output g29219;
output g29220;
output g29221;
output g30327;
output g30329;
output g30330;
output g30331;
output g30332;
output g31521;
output g31656;
output g31665;
output g31793;
output g31860;
output g31861;
output g31862;
output g31863;
output g32185;
output g32429;
output g32454;
output g32975;
output g33079;
output g33435;
output g33533;
output g33636;
output g33659;
output g33874;
output g33894;
output g33935;
output g33945;
output g33946;
output g33947;
output g33948;
output g33949;
output g33950;
output g33959;
output g34201;
output g34221;
output g34232;
output g34233;
output g34234;
output g34235;
output g34236;
output g34237;
output g34238;
output g34239;
output g34240;
output g34383;
output g34425;
output g34435;
output g34436;
output g34437;
output g34597;
output g34788;
output g34839;
output g34913;
output g34915;
output g34917;
output g34919;
output g34921;
output g34923;
output g34925;
output g34927;
output g34956;
output g34972;
output g24168;
output g24178;
output g12833;
output g24174;
output g24181;
output g24172;
output g24161;
output g24177;
output g24171;
output g24163;
output g24170;
output g24185;
output g24164;
output g24173;
output g24162;
output g24179;
output g24180;
output g24175;
output g24183;
output g24166;
output g24176;
output g24184;
output g24169;
output g24182;
output g24165;
output g24167;

wire 	g5057,g2771,g1882,g6462,g2299,g4040,g2547,g559
	,g640,g3017,g3243,g452,g464,g3542,g5232,g5813
	,g2907,g1744,g5909,g1802,g3554,g6219,g807,g6031
	,g6027,g847,g976,g4172,g4372,g3512,g749,g3490
	,g6005,g4235,g4232,g1600,g1714,g3649,g3625,g3155
	,g3355,g2236,g4555,g4571,g3698,g6073,g1736,g1968
	,g4621,g5607,g2657,g5659,g490,g311,g6069,g772
	,g5587,g6177,g6377,g6373,g3167,g5615,g4567,g3057
	,g3457,g6287,g1500,g2563,g4776,g4593,g6199,g2295
	,g1384,g1339,g5180,g2844,g1024,g5591,g3598,g4264
	,g767,g5853,g3321,g3317,g2089,g4933,g4521,g5507
	,g3618,g6291,g294,g5559,g5794,g6144,g3813,g562
	,g608,g1205,g3909,g6259,g5905,g921,g2955,g203
	,g6088,g1099,g4878,g5204,g5630,g5623,g3606,g1926
	,g6215,g3586,g291,g4674,g3570,g637,g5969,g6012
	,g1862,g676,g843,g4132,g4332,g4153,g5666,g5637
	,g6336,g622,g3506,g4558,g6065,g6322,g6315,g3111
	,g117,g2837,g939,g278,g4492,g4864,g1036,g128
	,g1178,g3239,g718,g6195,g1135,g6137,g6395,g3380
	,g5343,g554,g496,g3853,g5134,g1422,g1418,g3794
	,g2485,g925,g48,g5555,g878,g875,g1798,g4076
	,g2941,g3905,g763,g6255,g4375,g4871,g4722,g590
	,g6692,g6668,g1632,g5313,g3100,g3092,g1495,g6497
	,g6490,g1437,g6154,g1579,g1576,g5567,g1752,g1917
	,g744,g3040,g4737,g4809,g6267,g3440,g3969,g4012
	,g1442,g5965,g4477,g1233,g4643,g5264,g6329,g6351
	,g2610,g5160,g5360,g5933,g1454,g753,g1296,g3151
	,g2980,g6727,g3530,g4742,g4104,g1532,g4304,g2177
	,g3010,g52,g4754,g1189,g2287,g4273,g1389,g1706
	,g5835,g1171,g4269,g2399,g3372,g4983,g5611,g3661
	,g4572,g3143,g2898,g3343,g3235,g4543,g3566,g4534
	,g4961,g6398,g4927,g2259,g2819,g4414,g5802,g2852
	,g417,g681,g437,g351,g5901,g2886,g3494,g5511
	,g3518,g1604,g4135,g5092,g4831,g4382,g6386,g479
	,g3965,g4749,g2008,g736,g802,g3933,g222,g3050
	,g5736,g1052,g58,g2122,g2465,g6483,g5889,g4495
	,g365,g4653,g3179,g1728,g2433,g3835,g6187,g4917
	,g1070,g822,g6023,g914,g5339,g5335,g4164,g969
	,g2807,g5424,g4054,g6191,g5077,g5523,g3680,g3676
	,g6637,g174,g1682,g355,g1087,g1083,g1105,g2342
	,g6307,g3802,g6159,g2255,g2815,g911,g43,g3983
	,g1748,g5551,g5742,g3558,g5499,g2960,g3901,g4888
	,g6251,g6358,g1373,g157,g2783,g4281,g4277,g3574
	,g2112,g1283,g433,g4297,g4294,g5983,g1459,g1399
	,g758,g5712,g4138,g4639,g6537,g5543,g1582,g3736
	,g5961,g6243,g632,g1227,g3889,g3476,g1664,g1246
	,g6128,g6629,g246,g4049,g4449,g2932,g4575,g4098
	,g4498,g528,g5436,g16,g3139,g102,g4584,g142
	,g5331,g5831,g239,g1216,g2848,g5805,g5798,g5022
	,g4019,g4000,g1030,g3672,g3668,g3231,g1430,g1426
	,g4452,g4446,g2241,g1564,g6148,g6140,g6649,g110
	,g884,g881,g3742,g225,g4486,g4504,g5873,g5037
	,g2319,g5495,g4185,g5208,g2152,g5579,g5869,g5719
	,g1589,g5752,g6279,g5917,g2975,g6167,g4005,g2599
	,g1448,g3712,g2370,g5164,g1333,g153,g6549,g4087
	,g4801,g2984,g3961,g5770,g962,g101,g4226,g4222
	,g6625,g51,g1018,g4045,g1467,g2461,g5706,g457
	,g2756,g5990,g471,g1256,g5029,g6519,g4169,g1816
	,g4369,g3436,g5787,g4578,g4459,g3831,g2514,g3288
	,g2403,g2145,g1700,g513,g2841,g5297,g3805,g3798
	,g2763,g4793,g952,g1263,g1950,g5138,g2307,g5109
	,g5101,g5791,g4664,g2223,g5808,g6645,g2016,g5759
	,g3873,g3632,g3654,g2315,g2811,g5957,g2047,g3869
	,g3719,g5575,g46,g3752,g3917,g4188,g4191,g1585
	,g1570,g4388,g6275,g6311,g4216,g4213,g1041,g2595
	,g2537,g136,g4430,g4564,g3454,g3447,g4826,g6239
	,g3770,g232,g5268,g6545,g2417,g1772,g4741,g5052
	,g5452,g1890,g2629,g572,g2130,g4108,g4308,g475
	,g990,g1239,g31,g3412,g45,g799,g3706,g3990
	,g5385,g5881,g1992,g3029,g3171,g3787,g812,g832
	,g5897,g4165,g3281,g3303,g4455,g2902,g333,g168
	,g2823,g3684,g3639,g5327,g3338,g5406,g3791,g269
	,g401,g6040,g441,g5105,g3808,g9,g3759,g4467
	,g3957,g4093,g1760,g6151,g160,g5445,g5373,g2279
	,g3498,g586,g869,g859,g2619,g1183,g1608,g4197
	,g4194,g5283,g5276,g1779,g2652,g5459,g2193,g2393
	,g5767,g661,g4950,g5535,g2834,g1361,g3419,g6235
	,g1146,g2625,g150,g1696,g6555,g3385,g3881,g6621
	,g3470,g3897,g518,g3025,g538,g2606,g1472,g6113
	,g542,g5188,g5689,g1116,g1056,g405,g5216,g6494
	,g6486,g4669,g5428,g996,g4531,g2860,g4743,g6593
	,g2710,g215,g4411,g1413,g4474,g5308,g6641,g3045
	,g6,g1936,g55,g504,g2587,g4480,g2311,g3602
	,g5571,g3578,g468,g5448,g3767,g5827,g3582,g6271
	,g4688,g5774,g2380,g5196,g5396,g3227,g2020,g3976
	,g1079,g1075,g6541,g3203,g1668,g4760,g262,g1840
	,g70,g5467,g460,g6209,g74,g5290,g655,g3502
	,g2204,g5256,g4608,g794,g4023,g4423,g4537,g3689
	,g5381,g5685,g5681,g703,g5421,g862,g3247,g2040
	,g4999,g4146,g4633,g1157,g5723,g4732,g5817,g2151
	,g2351,g2648,g6736,g4944,g4072,g344,g4443,g3466
	,g4116,g5041,g5441,g4434,g3827,g6500,g5673,g5654
	,g3133,g3333,g979,g4681,g298,g3774,g2667,g3396
	,g4210,g4207,g1894,g2988,g3538,g301,g341,g827
	,g6077,g2555,g5011,g199,g6523,g1526,g4601,g854
	,g1484,g4922,g5080,g5863,g4581,g3021,g2518,g2567
	,g568,g3263,g6613,g6044,g6444,g2965,g5857,g1616
	,g890,g5976,g3562,g1404,g3723,g3817,g93,g4501
	,g287,g2724,g4704,g22,g2878,g5220,g617,g316
	,g1277,g6513,g336,g2882,g933,g1906,g305,g8
	,g3368,g2799,g887,g4912,g4157,g2541,g2153,g550
	,g255,g1945,g5240,g1478,g3080,g3863,g1959,g3480
	,g6653,g6719,g6715,g2864,g4894,g5677,g3857,g499
	,g5413,g1002,g776,g28,g1236,g4646,g2476,g1657
	,g2375,g63,g358,g896,g967,g3423,g283,g3161
	,g2384,g3361,g6675,g6697,g4616,g4561,g2024,g3451
	,g3443,g2795,g613,g4527,g1844,g5937,g4546,g3103
	,g3096,g2523,g2643,g6109,g1489,g5390,g194,g2551
	,g5156,g3072,g1242,g47,g1955,g6049,g3034,g2273
	,g6711,g4771,g6098,g3147,g3347,g2269,g191,g2712
	,g626,g2729,g5357,g4991,g6019,g6000,g4709,g6419
	,g6052,g2927,g4340,g5929,g4907,g3298,g4035,g2946
	,g918,g4082,g2036,g577,g1620,g2831,g667,g930
	,g3937,g5782,g817,g1249,g837,g599,g5475,g739
	,g5949,g6682,g6105,g904,g2873,g1854,g5084,g5603
	,g4219,g2495,g2437,g2102,g2208,g2579,g4064,g4899
	,g2719,g4785,g5583,g781,g6173,g6369,g2917,g686
	,g1252,g671,g2265,g6283,g6365,g5320,g6459,g901
	,g5527,g4489,g1974,g1270,g4966,g6415,g6227,g3929
	,g5503,g4242,g5925,g1124,g4955,g5224,g2012,g6203
	,g5120,g2389,g4438,g2429,g2787,g1287,g2675,g66
	,g4836,g1199,g5547,g3782,g6428,g2138,g2338,g4229
	,g6247,g2791,g3949,g1291,g5945,g5244,g2759,g6741
	,g785,g1259,g3484,g209,g6609,g5517,g2449,g2575
	,g65,g2715,g936,g2098,g4462,g604,g6589,g1886
	,g6466,g6346,g429,g1870,g4249,g6455,g3004,g1825
	,g6133,g1008,g4392,g5002,g3546,g5236,g1768,g4854
	,g3925,g6509,g732,g2504,g1322,g4520,g2185,g37
	,g4031,g4027,g2070,g4812,g6093,g968,g4176,g4405
	,g4408,g872,g6181,g6381,g4765,g5563,g1395,g1913
	,g2331,g6263,g50,g3945,g347,g5731,g4473,g1266
	,g5489,g714,g2748,g5471,g4540,g6723,g6605,g2445
	,g2173,g4287,g2491,g4849,g2169,g2283,g6585,g121
	,g2407,g2868,g2767,g1783,g3310,g1312,g5212,g4245
	,g645,g4291,g79,g182,g1129,g2227,g6058,g4204
	,g2246,g1830,g3590,g392,g1592,g6505,g6411,g1221
	,g5921,g106,g146,g218,g6474,g1932,g1624,g5062
	,g5462,g2689,g6573,g1677,g2028,g2671,g34,g1848
	,g3089,g3731,g86,g5485,g2741,g2638,g4122,g4322
	,g5941,g2108,g25,g1644,g595,g2217,g1319,g2066
	,g1152,g5252,g2165,g2571,g5176,g391,g5005,g2711
	,g1211,g2827,g6423,g4859,g424,g1274,g85,g2803
	,g6451,g1821,g2509,g5073,g1280,g4815,g6633,g5124
	,g6303,g5069,g2994,g650,g1636,g3921,g2093,g6732
	,g1306,g5377,g1061,g3462,g2181,g956,g1756,g5849
	,g4112,g2685,g2197,g6116,g2421,g1046,g482,g4401
	,g6434,g1514,g329,g6565,g2950,g4129,g1345,g6533
	,g3274,g3085,g4727,g1536,g3941,g370,g5694,g1858
	,g446,g4932,g3219,g1811,g3431,g6601,g3376,g2441
	,g1874,g4349,g6581,g6597,g5008,g3610,g2890,g1978
	,g1612,g112,g2856,g6479,g1982,g6661,g5228,g4119
	,g6390,g1542,g4258,g4818,g5033,g4717,g1554,g3849
	,g6704,g3199,g5845,g4975,g790,g5913,g1902,g6163
	,g4125,g4821,g4939,g3207,g4483,g3259,g5142,g5248
	,g2126,g3694,g5481,g1964,g5097,g3215,g111,g4427
	,g7,g2779,g4200,g1720,g1367,g5112,g19,g4145
	,g2161,g376,g2361,g582,g2051,g1193,g5401,g3408
	,g2327,g907,g947,g1834,g3594,g2999,g5727,g2303
	,g3065,g699,g723,g5703,g546,g2472,g5953,g6439
	,g1740,g3550,g3845,g2116,g3195,g3913,g1687,g2681
	,g2533,g324,g2697,g5747,g4417,g6561,g1141,g2413
	,g1710,g6527,g6404,g3255,g1691,g2936,g5644,g5152
	,g5352,g6120,g2775,g2922,g1111,g5893,g1311,g3267
	,g6617,g2060,g4512,g5599,g3401,g4366,g94,g3129
	,g3329,g3325,g5170,g4456,g5821,g6299,g3727,g2079
	,g4698,g3703,g1559,g943,g411,g3953,g3068,g2704
	,g6035,g6082,g49,g1300,g4057,g5200,g4843,g5046
	,g2250,g319,g4549,g2453,g5841,g5763,g3747,g2912
	,g2357,g164,g4253,g5016,g3119,g1351,g1648,g4519
	,g5115,g3352,g6657,g4552,g3893,g3211,g929,g5595
	,g3614,g2894,g3125,g3821,g4141,g4570,g5272,g2735
	,g728,g6295,g5417,g2661,g1988,g5128,g1548,g3106
	,g4659,g4358,g1792,g2084,g3061,g3187,g4311,g2583
	,g3003,g1094,g3841,g4284,g3763,g3191,g4239,g3391
	,g4180,g691,g534,g5366,g385,g2004,g2527,g5456
	,g4420,g5148,g4507,g5348,g3223,g4931,g2970,g5698
	,g3416,g5260,g1521,g3522,g3115,g3251,g1,g4628
	,g1996,g4515,g4300,g1724,g1379,g12,g1878,g5619
	,g71,g59,g7266,I11691,I13054,I13149,I13152,I13031
	,I12994,I13010,I13020,I13252,I12991,I12935,g9901,g10108
	,g7231,g9688,g9964,g9820,g8286,g10030,g9819,g8456
	,g9581,g10176,g8571,g9902,g8356,g9689,g9822,g9748
	,g10073,g9636,g9821,g10109,g9534,g9965,g9332,g9686
	,I14827,I14679,I14970,I14742,I15073,I14902,I14797,I15030
	,I14866,I14905,I14839,I14241,I14935,I14301,I15162,I14773
	,I14271,I14893,I14999,I14222,I14896,I14967,I14836,I14079
	,I15070,I14932,g8989,g9153,g9637,g9213,g9186,g9154
	,g9245,g9478,g9477,g9280,g6869,I13847,g9716,g8579
	,g9590,g9629,g9574,g7379,g8626,I12666,g10154,g9480
	,g9049,I12963,g9056,g7251,I13109,g8530,g9413,g9640
	,g7356,g10341,g9518,g7850,I12135,g8899,I18700,g9246
	,g9086,g10274,g6818,g7673,I12861,g6958,g8021,g8770
	,I12109,g8218,g10185,g7395,I15190,I12840,I12902,I12899
	,g9250,g9970,I16606,I17852,g9916,g7964,g9177,g9060
	,g10261,g8733,g9456,g9283,g10199,g7785,g10205,g10160
	,I15144,g7344,g6804,g7537,g7297,I12016,g8859,g9959
	,I18734,g8011,I13723,g8479,I12372,g8068,g8632,I12611
	,g10034,g9968,g7947,I12314,g8138,g7557,g7535,g9490
	,g8131,g7928,I11824,g7227,g7163,g7072,g9339,I12096
	,g7778,g10266,g9300,g7518,g8967,g8914,g8830,I12003
	,g7049,I16168,I18066,I13509,g6994,g8234,g7235,g7162
	,g7026,g8728,g9713,I17819,g8458,I13240,g9618,g9742
	,I13317,I12401,I12061,g10032,I12159,g8945,g7661,g7918
	,g9174,g7851,g7696,g6800,g9397,g7868,g9664,g7846
	,g7991,g7840,g7521,I18555,I18509,g7470,g9591,g8302
	,g9462,I12199,g8575,g9602,g7788,I15208,g7496,I18560
	,I18728,g7471,g9694,g7322,g8898,g9220,g7655,I12927
	,g9985,g7932,g7437,I18694,I16795,g7394,g10050,g7087
	,g9162,I12086,g7985,g7132,g7187,g7563,I18662,g10207
	,g7513,I18614,I12344,I13694,I11685,g10084,g7404,g8608
	,g10222,I11753,g7809,g7548,g9663,g8803,g7017,I13684
	,g9967,g7715,g10074,g10002,I12203,g7069,I11801,g10169
	,g8155,I13360,g9856,g6808,I12144,g8951,g6803,g6926
	,g9671,g9011,I18337,I18297,g8955,I12523,g8345,g9654
	,g8373,g7301,I12415,I16328,I16417,g8904,g7666,g8690
	,g8681,I11992,g7685,g7495,g7259,g8889,g9852,g7828
	,I12013,g8851,I15732,g7591,I18709,g10043,g10124,g7296
	,I15102,g8438,g8216,I12451,g7876,g10058,I13374,g9818
	,I12217,I13139,g9460,g8091,I13892,g9639,g8249,I12089
	,g8745,g7975,g8673,g8133,I12411,g6900,g8751,g9771
	,I17857,I17999,g9714,g7886,g10159,I13875,g7285,I16847
	,g7472,I15238,g7439,g8381,g7002,g7167,g7138,I12261
	,g7619,g6873,I13581,g10102,g8906,g8165,g6990,g7670
	,I13065,g9252,I13037,g9648,g9015,g8388,I12336,g6987
	,g9700,g7335,g9018,I11726,g6830,g8002,g9691,g9510
	,g7304,g8609,g8407,g8964,g9832,g9360,g8177,g9064
	,g9661,I17964,I12735,g8217,g6874,g8663,I13729,g7228
	,g7191,g8715,g10180,g8686,I11903,g7258,g9887,g9333
	,g9903,I12997,g7834,g8281,g6904,g9239,g8070,I13744
	,g7267,g9724,g9669,g8847,g9775,g7063,g7469,g7289
	,g10191,g7410,g8836,g9905,I14563,g8679,g9092,g8340
	,g9733,g7913,I12538,g10152,g7424,g7092,g8720,g8721
	,I12719,g7836,g7690,g8606,g8864,g8107,g7275,g7423
	,g8228,g9620,g6820,g7750,g7777,g7216,I16770,g7443
	,I18600,I11701,g9483,g7903,g8639,g9442,g9379,g8700
	,I11716,g9684,g7073,g9989,I12176,g9311,I17938,g8086
	,g9969,g7499,g9050,g8654,g9007,I18333,I12240,g8267
	,g8565,g8659,g7400,I11860,I16246,g9662,g9537,g9316
	,g9557,g7027,g7763,g6991,g7497,I18752,g7582,g8033
	,g8635,I12848,g8840,I12819,g9973,g7450,g10123,I13623
	,g7438,I16821,I15837,g8301,I19837,I12123,g8651,g7158
	,g9807,g6954,g7202,g7096,g9745,I12608,g8443,g9217
	,g6814,I12120,g9000,I12577,I15536,g8442,g8863,I11655
	,g8056,g9954,g9889,I13382,g8296,g8756,g7261,I11908
	,g7764,g6957,I12749,g6989,g7636,I12805,I12360,g8046
	,g9800,g9730,I11632,g10106,g8154,I13637,I13749,g10275
	,g8297,I16713,g9888,I13442,g8363,g9223,g9932,g9681
	,I13276,g10338,g9670,I18107,I16639,g7549,I16181,I18092
	,g7948,g8685,g9091,g9051,I18360,g7293,I11896,g7246
	,g10038,g7675,g9226,g9958,I13280,g9683,I13287,I16357
	,I16345,g8075,g8457,g10184,g10312,g9451,g9253,g9595
	,g8211,g9500,I14619,g6846,g9392,I12189,g7170,I11665
	,g8092,g7184,g9739,g7804,g9816,I14424,g9601,g7462
	,g9100,g8507,g9206,g7601,g8240,g7995,g9407,I12746
	,g7697,g7892,g9509,g9449,g7517,I11835,I12893,I12903
	,I12837,I12572,g8734,I12277,g10158,g7157,I11682,g9978
	,g9992,g7064,g7446,g7134,g9962,g7824,g10036,g8497
	,g9880,g6997,I12793,g10308,g8566,I13518,g8531,g6895
	,g9913,g7511,g6841,g10150,g9158,g10119,g9853,g7018
	,g8592,I12563,g8399,g9657,g9030,g7597,g7577,g10079
	,g9729,g9594,g9728,I13166,g9498,g7046,g8650,g8905
	,g9390,g9644,g9933,g8958,g8172,g9600,I16217,g9552
	,I14395,g9760,g9012,g8125,I11820,g9180,I12355,g9203
	,g8449,I12782,I12761,I14450,I12654,g8364,I12605,I15542
	,I11877,I12887,I12884,g10183,g9976,I13708,g10139,g7149
	,I11743,g8539,g8343,I12519,g8764,g8713,g7086,g8227
	,g8170,I13497,g8406,g7095,g10153,g6848,g7315,g9229
	,g9616,I13236,g9753,g9835,g7490,I12103,g8766,g7680
	,g7567,I12583,g8186,I12580,g10197,I11626,g8538,I12333
	,I15036,g9099,g8623,g6941,g9434,g9511,g6840,g10151
	,g8097,g8059,g8558,g7197,g9334,g7118,g7765,g8691
	,g9551,I16193,I14365,g9496,g6917,g6918,g8584,I18795
	,I12618,g8534,g7139,g9678,g6923,g8136,g10166,g7396
	,I13202,g9554,g8123,g10072,I11635,g8593,I11737,I12758
	,g7733,g9538,g8146,g10000,g8287,g7023,g7153,g10081
	,g8541,I12117,g10262,I16401,I16391,g9705,g8418,g8462
	,g9337,I12767,I12764,g7512,I18504,g7436,I18460,I13564
	,g10040,g9861,g10086,g10203,g10096,g10110,g10281,g9444
	,g9152,g8163,g8112,g7845,g9055,g9073,g10179,g9472
	,g8390,g8229,g8397,g9187,g8005,g9535,g10136,g9374
	,I13424,g9927,I15824,I19818,g8239,g8182,I12468,g8037
	,g10026,g9744,I13321,g8672,g6985,g9439,g9070,I12074
	,g9906,g7749,g6982,g6986,g8292,I12503,g7232,g6831
	,g7779,I11750,I15663,g8426,g9900,g7405,I12418,g9077
	,g8330,g9699,g6802,g9556,I13206,g8669,g9808,g7970
	,g7827,g9883,g9103,g9506,I13462,g9264,g9754,I17901
	,g9982,I18293,g8954,g8903,I18276,g10060,g9586,g7308
	,g8180,g9752,I11688,I13077,g9402,I13606,g7631,g7343
	,I16762,g10033,g6903,g7236,g7183,g8833,I12112,I16201
	,I13726,I12644,g8587,g9305,I18653,g9582,g10047,g7441
	,g7411,I12437,g8179,I13352,g7963,g10311,g7532,g7917
	,I12300,g7519,g8087,g7262,g9450,g8316,g10229,g6995
	,g7684,g7541,I12026,g7340,g8113,g9364,g9797,I11864
	,g8508,I13182,g9527,I18813,I15677,g8106,g8718,g8765
	,g6887,g6825,g7806,g8522,g8561,g7952,g8224,g9977
	,g8492,I12783,I12779,I12776,g8201,g8461,g6809,g9194
	,g9559,g7431,g9715,g8829,g7109,g6799,g10027,g7352
	,g8526,g7224,I12287,g9372,g9298,g9321,I13699,g9291
	,g9974,g7461,g10143,I12083,g10190,g7192,g9898,g9274
	,g9585,g7442,I13718,g7397,g7536,I18609,g7960,g9429
	,g8171,I11816,g8519,I13094,g9839,g10318,g7116,g7780
	,g9214,I12064,g6827,g9899,g7564,g6816,g7362,g9479
	,g7523,g10028,g9095,I16371,g7908,I13473,g6953,g10118
	,g9649,g7280,g8743,g8237,g8434,g8387,g8080,I13452
	,g9907,g8505,I18758,I16829,I16741,g8026,g9040,g9862
	,g7635,g8748,I12033,g10175,I11623,g8055,g8350,g8324
	,g9485,g8187,g10082,I13705,g8678,g8806,g8848,g7475
	,g8500,g7926,g8160,g8631,g7980,g9911,g9061,g8441
	,g10224,I16875,g7498,I15284,g7473,g6978,g10223,g9828
	,g8504,I12487,g8280,g8854,I12046,g10232,g9826,g8478
	,g8278,I12483,g10155,g9999,g7867,g9672,I12544,g8362
	,I12541,g10181,g6849,g9779,g8105,g8102,g7907,g8300
	,I12631,I12382,g10133,I11793,g8334,g10039,I18845,g7175
	,g7209,g9815,g8480,g8696,g9831,I12106,g9083,g9491
	,I13124,I11777,g10044,g7898,I18825,I15697,g8933,g8883
	,g6984,g9523,g7174,g8643,g8347,I12790,I12910,I12858
	,I12811,g8928,I16575,g6940,g8742,g8804,g7544,g8567
	,g10157,g8997,I12132,g9638,g9071,g7528,g9806,g10320
	,g7863,g9166,I12141,g8895,g9679,I12067,g8725,g7110
	,g10099,g10001,g7841,g10078,g9369,g9036,I12890,g9762
	,g7456,g9546,g10217,g8205,g9834,g7781,g7611,g7927
	,g7650,g8984,g6992,g8938,I12183,g9354,g8796,g8774
	,I12049,g9891,I16803,g8583,g8680,g7957,g8858,g9759
	,I18835,g7393,I18647,g10172,g9381,g10206,g9827,g7349
	,g7953,g7345,g9569,g9863,g9984,g6956,I12251,g6996
	,g9541,g9326,I13043,g7392,g9416,g8655,g10156,I11980
	,I13326,g8400,g7716,g8506,g9892,g10200,g8957,I12896
	,g7880,g9492,I11809,g10194,I12070,g8948,g7487,g8164
	,g9269,g9833,g9704,I13007,I12172,g9285,g7909,g9848
	,I12151,g9044,g9693,g10022,g9212,g9626,I15717,g9338
	,g10057,g9014,I13390,g9824,g9951,g7479,g7178,I12493
	,g8284,g10085,g8677,g9575,g9690,g6836,g9543,g8150
	,g8607,I17970,g9755,g7451,I12463,g8236,g9946,g6837
	,g7219,I11892,g7244,g9568,I13539,g10053,g6988,g7943
	,g8956,g7380,I12534,g7592,g9501,I11734,g7873,g9443
	,g8769,g6811,g9766,I12056,g9380,g9761,g9542,I12728
	,I12950,g9020,g9013,g7701,g7693,g9415,g6847,g10115
	,I13552,g10083,g8195,I17932,g9599,g9536,g7922,I13634
	,g8807,g7374,g9890,I12773,I13401,g7998,g7252,g7212
	,g9197,I13672,g8990,g8290,g6826,g9960,g8093,g7150
	,g9613,g9309,g7520,g7142,g9631,g9645,g8255,g10042
	,I12227,g10037,g6870,g8219,g6999,I13329,g9805,g9708
	,I12041,g7643,g9920,I12907,I12808,g9910,g7195,g8808
	,I12030,g8259,g6829,g10289,g7854,g7327,g9598,I12167
	,g9259,g6801,g8404,I12568,g6855,g8052,g9621,g6993
	,g8714,g8181,g7553,I13740,g8616,g10059,g10117,g9776
	,g7939,g8354,I12530,g9299,g9778,g9072,g7891,g7268
	,g9971,g10213,g7533,g7247,g7936,g9698,I12269,g6817
	,g9692,g9934,g10204,g6854,g7328,g9567,g9516,g7387
	,g7972,g6819,g8183,g9467,g8466,g7440,g9576,g7649
	,g9685,g9842,I17814,g8431,g7888,g8944,g10130,g10111
	,g6839,g6998,g8440,g8064,g9653,g7361,g10290,g8977
	,I12930,I12826,g7992,g9909,g9484,I13057,g10019,g10080
	,I18667,g7522,g10212,g7752,g8872,g8514,g7971,g7239
	,g8088,g8594,g7514,I18778,g7050,g9619,g8822,I12092
	,g9003,g10120,g9517,g7835,g7040,g8741,g8676,g10335
	,g9373,g10178,g6845,g8697,g9732,g9721,I11843,g7222
	,g9963,I12876,I12770,g10035,g7534,g9777,I11629,g10140
	,I11721,g9284,g8890,g7418,I12000,g8891,g8310,g7870
	,g9792,g8540,g10121,g7933,g7858,g10177,g9386,g9489
	,g8620,g6810,g9282,I11785,g10093,g10014,g7314,g8346
	,g6927,g10114,I13334,g10182,g9914,g7802,g10219,g9875
	,I13597,I12214,g9529,g10116,g9751,g9630,g9961,g9749
	,g9924,g7041,g7003,g9499,g10129,g9564,g9184,g8612
	,I17787,g9660,g8365,g8396,g7805,I13548,g8439,I17892
	,g9234,g9740,g8119,g6983,g8666,I11708,g9247,g8137
	,g8057,g6850,g9995,I13483,g9809,I12497,g6828,g8451
	,g8630,g9607,g9829,g8273,g9558,g9931,g8553,g9037
	,I12128,g10337,g8341,g7503,g8139,I11740,g9257,I11697
	,g8644,g6815,g8389,g8450,g8509,I11746,g9547,g10147
	,g9860,g10231,g10112,g9614,g9200,g8009,g7686,g9024
	,I12954,g8241,g10113,g8477,I12855,g7166,g7627,I12823
	,g9843,I12787,g9915,g8282,I12709,g8591,g9983,g8016
	,g8912,g8744,g9731,g8993,g9414,g10218,g9804,g6959
	,g10334,g9433,g6975,g10090,g10165,g8647,g7751,g8114
	,g8058,I11617,I11620,g6960,g10278,g7369,g8130,g10077
	,g6838,g7581,I12987,g7115,g9488,I13715,I12799,I12712
	,g10430,g10364,g12076,g12180,g12181,g12036,g11964,g11984
	,g12012,g12321,g11963,g11912,g12074,g12217,g10877,g11988
	,g12109,g12038,g11165,g12143,g12037,g11204,g11949,g12322
	,g11235,g12075,g11182,g11989,g12041,g12013,g12182,g11965
	,g12040,g12218,g11928,g12110,g11867,g11985,g8712,g8805
	,g10287,g10520,g9104,g11869,g10603,g10585,g10380,g6755
	,g6754,g11618,g11527,g11483,g12220,g12294,I15128,I14609
	,g10537,I13995,I14033,I12878,g11414,g11360,g8703,I12204
	,g8791,g10820,g8841,g12797,g11018,g8876,g11345,g11273
	,g12117,g12114,g11953,g12079,g9021,g10614,g12687,g12762
	,g11006,I12345,g11171,g10921,I14712,I15174,g12296,g12201
	,g11708,g6974,g10808,g10998,g10841,g10677,I14204,g11382
	,g6875,I13044,g6972,g11934,g12016,g11914,g12113,g12817
	,g11366,g7640,I24033,I24054,g12346,g12249,g12194,g12225
	,g12023,g12483,I13403,g10884,g10626,g10922,g11003,I12289
	,g8285,g9935,g12252,g12830,g11126,g10362,g10684,g6905
	,g11412,g10388,g11010,g12292,I14764,g12235,g12646,g12553
	,g11205,g10029,g12190,g11994,g12148,g11441,I12241,g11046
	,g12027,g12344,g10401,I13336,g10598,I14991,I12270,g12752
	,g10581,g7812,g10087,I24530,I24552,g10759,I15333,g11244
	,g11954,I24603,I24585,g7028,I15041,g11384,I24508,I24527
	,g11330,g12116,g7515,g10586,g11939,I14350,g11607,g6946
	,I14505,g6772,I12877,I14050,g7161,g12160,g11027,g10622
	,g12228,g10403,I14267,g11201,g7618,g11834,g11804,g12099
	,g12476,g10556,g10827,g12358,g11127,g9281,g10617,g10573
	,g8844,g8974,g11972,g10625,g10609,I14508,g11374,g11270
	,g10654,g12043,g12680,g12632,g10715,g10699,I11866,g10356
	,g10760,g10587,g10568,g11996,g10653,I12271,I12374,g12526
	,I13511,g10550,g11969,g10615,g12234,g12126,g12163,g12121
	,I13391,g12466,g12318,g10319,g10565,g11148,g12550,g10489
	,g7704,g11958,g11017,g11957,g12118,g12083,g7542,g8818
	,g8922,g12399,g7558,g12289,I14567,g12065,g9747,g10398
	,g10367,I15253,g7831,g11995,g12082,g10428,I13078,g11862
	,g12078,g11952,g11047,g10198,g10934,g11130,g11945,I13184
	,g10529,g11216,I12470,g10578,I12253,g10141,I12729,g11469
	,g12795,g11355,g12045,g10031,g10611,g11012,g10862,g12088
	,g12486,I12730,g7586,I14584,g10354,I14883,g6961,g10799
	,g8355,g12022,g12435,g10391,g12314,g10427,g10003,g11142
	,I14955,I13862,I24582,I24555,g10602,g11956,I14326,g12149
	,g12021,g12374,g10360,I14247,I12098,g12794,g12308,g11115
	,g10873,g12361,g12523,g11911,g7674,g7717,g9185,g12695
	,g12297,g12604,g10665,I14275,g7596,g7097,g10656,g9746
	,g7474,g10683,g12419,g12780,g10519,g12744,g10387,I12252
	,g10349,g12622,g12831,g10421,g11173,g11232,g12601,g12505
	,g12453,g12244,g11380,g7566,g11797,g11773,g7753,g11034
	,g10604,g11960,g11023,g12418,g12256,g10413,g7595,g7659
	,g11950,g11913,g11968,g11933,g11029,I15382,g7647,g10377
	,g10664,g8821,g8879,g8925,g8792,g11449,g12461,g11283
	,g11203,g7004,g9417,g7624,g11940,I12545,g11924,g12417
	,I15262,g7051,g12416,I13453,g8085,g8515,I14381,g10624
	,g10623,g10971,g10946,g12311,g12154,g11172,g7565,g11279
	,g12821,g12822,g10383,g12364,g11948,g11881,g11383,I13464
	,g11653,g11346,g11566,g11303,g11033,g10601,I14158,g10272
	,g12085,g11935,g11991,g11998,g11977,g12226,g6756,I14475
	,g7543,g11846,g12015,g12170,g11020,g11715,g11415,g11833
	,g11697,g11223,g11026,I12219,I13498,g12050,I15340,g10379
	,g9917,g11107,I14054,g10796,g10584,g12019,g10355,I14816
	,g10358,g7594,g10582,g10416,g9340,g7117,g10755,g12415
	,g10288,g10632,g12739,g12347,g10490,g12700,g12465,g7615
	,g12025,I13520,g10233,I12288,g10970,I11826,g12179,g10415
	,g10605,g12147,g11993,g12188,g12432,g8790,I24030,I24018
	,g11357,g11043,g10357,g10726,I12076,g10368,I14257,g12413
	,I13183,I11865,g12198,g11035,I24524,I13937,g10395,I13565
	,g12151,g11975,g12119,g11117,g9772,g12014,g12042,g11309
	,g11753,g8542,g10724,I13731,g7626,I13750,g10555,g10374
	,g11741,I14480,g12197,g10107,I13079,g6868,I14225,I13443
	,g12017,g11445,I13463,g12246,g11866,g10831,g11396,g12196
	,g10351,g12227,g12053,g12287,g12540,g8135,I14046,I24003
	,I24015,g12341,g6976,g11030,g10389,g10386,I12075,g11028
	,g12317,I12469,g8417,g10909,g10905,g12204,g12804,g9864
	,g11114,g12443,g12738,g12772,I12279,g12812,I14185,g11584
	,g11754,g11763,g12467,g12806,g12755,g10951,I15250,g12779
	,I15087,g10695,g10649,g12024,g12195,g12122,g7632,g11885
	,g10402,g12018,g11245,I13979,g8778,g6971,g6789,I14550
	,I12402,I13383,g10376,g12295,g11276,g11735,g8481,g10706
	,g10371,g10373,g11042,g11563,g11473,g11435,g12571,g12805
	,g12824,g11446,g10375,g10898,g12185,g7993,g6767,I14455
	,g11812,g10881,g10872,g10621,I13066,g10674,g10719,g7623
	,g10610,g11978,I24546,g10566,g11992,g10618,g10370,I13499
	,g10411,g11190,g6973,I11879,I15205,g10273,I11878,g8470
	,I14409,g8572,g11119,g8032,g7121,g11666,g11884,I13110
	,g10406,g12125,g12081,g10800,g11200,g10397,I15223,I15002
	,g10361,g10366,I13519,g8795,g10396,g12046,I14119,g10405
	,I14593,g6856,g11427,g11544,g8405,g8921,I12841,g7148
	,g11231,g11261,I13968,g8757,g10541,g11134,g10897,g11849
	,g10652,g10882,g12823,g11413,I12263,g11907,I14862,g6832
	,g7766,g12659,g10540,g11976,g12051,g12192,g12437,g9687
	,g12255,g10966,g11149,g10980,g11513,g11786,g12233,g12008
	,I13751,g10142,I14537,g6782,g11841,g8038,g8812,I13990
	,g10392,g8763,g10381,g11889,I14823,g6821,g8411,g7633
	,g12768,g10795,g12345,g7634,g8476,g12307,I12850,I12849
	,g11815,g12428,g10393,g7196,I13141,g10960,g10917,g10518
	,g7738,g12135,g6928,g6888,g11892,g11999,g10551,g11714
	,g12054,g10708,g10414,g8357,g11039,g11083,g11679,g12464
	,g11496,g10407,g11811,g10323,g11861,g10420,g9155,I13730
	,g8740,g11493,g10856,g11031,g10359,g6955,g10893,g10390
	,g7994,g11344,g12284,g10918,g11736,g10497,g10061,g10369
	,g10400,g10961,g11363,g11122,g10372,g7617,g11971,g11955
	,g12189,I12218,g12073,g11251,g12166,g11865,g7526,g7502
	,g8134,g12086,g10378,g10353,g7660,g12778,g9780,g7074
	,g10410,I12205,g11721,g10216,g10399,g6977,g6867,g10230
	,I12346,g11927,g11385,g11692,g11796,g11658,g7616,g10409
	,g12245,I14570,g12440,g8971,g12369,g11214,g11779,g7791
	,g12708,g10564,g12047,g10725,g11810,g11233,g10350,g11472
	,g7689,g7593,g11110,g10404,g10394,I13510,g10408,g7516
	,g11316,I12097,g10412,I11825,g11038,I12373,g10295,g11832
	,g7527,g10352,g11888,g11762,g11910,g7625,g10382,g8880
	,g11011,g7648,g12259,g12323,g8595,g11769,I24505,I24482
	,g10736,I13111,g11915,g12581,g12111,g11951,g11621,I12842
	,I15212,g11443,g11411,g11610,g10883,I15078,g10511,g11320
	,g11967,g11252,g11191,g11213,g11155,g10510,g10803,g10821
	,g12405,g10822,g11489,g12207,g12035,I12403,g10896,I24616
	,g10929,g12232,g11426,g12343,g12459,g12115,g11674,g12124
	,g12521,g12356,g10567,g11932,g12306,g12588,g12463,g12587
	,g12159,g11707,g12186,g10878,I24051,g11044,g11312,g12152
	,g10829,g11546,g11639,g12589,g12525,I13140,g10528,g12080
	,I24048,g11543,g11424,g10501,g12357,g12288,g12153,g12000
	,g11397,I12262,g10802,g11163,g11747,I13067,g11858,g12219
	,g10569,g10793,I14923,g10666,g11248,g11394,g11442,g11497
	,I15051,g10928,g10709,g12651,g11019,I24579,I24597,g12052
	,g11326,g11729,I14289,g12761,g10616,I12242,g10890,g12193
	,g11959,g12084,g11395,g12340,g11016,g10935,g10939,g10561
	,I24067,I24075,g11037,I13384,g11024,I13444,g10515,g11491
	,g10947,I14198,g12515,g11997,I14788,g12087,g10967,g11903
	,g12593,g12785,I12278,g12522,g10675,g11045,g10704,g11184
	,g12412,g12208,g11537,g11356,g10801,g10819,g11979,g11306
	,I24549,I24027,g10707,g11891,g11302,g11490,g11961,g11313
	,g12371,g11970,g12145,g12293,g12411,I13566,I14516,g12798
	,g10916,I24064,g10999,g11937,g12591,g12169,g11036,I24576
	,g11893,g12711,g11990,g11740,g10583,g11002,I13850,g12048
	,I14228,g10676,I24600,g10671,g12662,g11675,g10552,g11370
	,g10948,g10619,g11669,I13454,g12120,g12729,g12044,g11676
	,g10655,g12429,I12546,g11755,g11409,g12527,I14733,g12639
	,I15121,g12150,g12049,g11938,g10899,g10657,g11780,I13045
	,I15363,I24619,I24625,g11116,I13392,g11974,I15306,g12146
	,g11936,g10902,g11916,I13402,g12333,g12112,g10720,g10732
	,g10705,g10491,g12479,g12020,g12222,g10925,g11381,g12460
	,g12730,I15298,g12638,I14853,g12223,g11973,g11280,I13335
	,I14169,g12847,g12850,g12848,g12855,g12856,g12852,g12846
	,g12854,g12849,g12853,g12851,I15587,I15533,I15650,I15556
	,I15705,I15623,I15569,I15682,I15609,I15626,I15593,I16452
	,I15636,I16535,I15736,I15564,I16486,I15617,I15667,I16438
	,I15620,I15647,I15590,I15448,I15702,I15633,g13494,g13412
	,g13302,g13087,g13070,g13051,g14562,g14357,g14198,g14173
	,I15474,I16521,I15788,I16613,I16135,I15906,I15577,I16555
	,I16476,I15782,I15915,I15893,I16460,I16709,I16498,I16057
	,I16090,I15929,I16040,I15600,I16117,I16479,I15773,I16502
	,I15550,I16102,I16077,I16526,I16150,g14415,g13081,g11631
	,I15341,g9391,g14361,g14940,g14902,g15036,g12578,g14861
	,g15008,g10874,g11562,g14178,g14254,g13336,g12885,g11571
	,g13955,g13920,g14094,g11470,I14276,I15193,I16671,g8871
	,g14313,g10733,g11514,g14008,g14041,g14234,g13959,g11533
	,g14335,I15147,g11372,g12835,g14408,g11293,g13913,g14011
	,g13980,g8069,g13291,g13006,g12982,g13464,g7133,g12909
	,g7620,g14758,g14953,g14656,g14915,g12402,g14879,g10823
	,g13540,g14124,g11269,g12905,g9972,g12887,g12901,g8124
	,g11401,g11677,g13662,g13756,g13727,g13511,g13527,g12839
	,g13326,g14874,I16646,g11123,g12950,g14943,g14864,g14587
	,g10553,g11691,g12101,g12628,g11160,g12173,g12902,g11429
	,g14048,g14075,g14151,g13923,g14192,g14248,I16695,g8010
	,I14964,g10365,g12891,I14939,I14481,g7803,g12904,g13541
	,g12749,g12497,I13857,g13492,g11609,g14165,g12838,g12871
	,I14713,g11181,g14097,g14218,g13806,g13831,g14002,g11250
	,g13155,g11291,g11178,g7823,g9461,I14249,g14612,g11430
	,g13872,g14028,g12865,g13059,g13288,I15241,g12897,g12941
	,g7879,g14177,g14182,g12866,g11025,g12721,g13567,g13986
	,g11480,g12692,g13322,g9295,g14417,g13627,g11129,g13834
	,g13345,g12883,g13314,g14589,g13265,g12843,I15003,g13868
	,I15088,g13628,g13486,g13469,g12546,g13954,g10307,g13000
	,g14061,g10608,g12558,g14848,g14885,g14051,g14018,g13941
	,g13909,g14596,g12899,g14867,g14232,g11236,I15334,g12908
	,g13566,I14510,g14101,g13873,g14098,g14069,g14566,I14956
	,g13911,g10828,g11702,g14851,g14807,g14438,g7857,g10542
	,g14392,g12886,g8873,g13273,g13315,g11170,g11512,g14407
	,g14545,g11510,g13121,g10741,g10761,I14186,g11981,g14030
	,g9823,g12879,g10504,g12884,g10678,g11192,g13973,g11592
	,I14258,I14833,g10336,g9904,g13570,I16143,g14506,g13699
	,g14004,g12107,g14148,g14126,g14892,g15018,g14858,g12512
	,g14968,g14810,g10869,g14614,I14884,g11771,g12944,g14895
	,g14813,g12009,g13708,g12492,g14755,g14841,g13134,g14981
	,g15014,g12716,g10627,g13739,g13634,g13995,g10429,g11249
	,g7887,g11724,g12067,g12577,g11139,g12129,g12898,I14817
	,g10981,g13035,g13493,g12889,g10533,g10738,g9975,g11194
	,g11479,g10721,g11217,g12859,I15004,g12381,g12002,g12449
	,g10588,g11111,g12059,g12890,g13432,g14418,g12900,g13523
	,g13330,g14446,g14170,g14082,g14058,g14142,g14021,g11534
	,g12735,I14398,g14237,g14085,g14024,g11143,g11448,g11398
	,g10762,g10794,g7223,I15033,g12367,g12903,g9966,g12862
	,g14792,g14644,g11467,g11450,g11128,g12867,g14999,g14855
	,g14933,g14735,g14127,g13889,g13892,g13915,g14208,g13048
	,I14368,g12864,g11207,g12863,g11444,g11238,g11519,g12869
	,g13080,g11166,g13795,g14816,g13794,g11640,g12645,g12767
	,g12796,I13802,g10658,g14586,g12896,g13507,g14212,I15263
	,g11509,g14202,g14190,g14680,I16618,g10041,g14752,g14665
	,g14959,g14927,g14956,g12430,g14791,g13729,g13595,g13569
	,g13624,g14868,g14822,g12915,g14825,g12945,g14157,g14055
	,g13963,g14116,I14187,g14918,g14627,g14723,g14800,g14659
	,g14683,g12563,g13103,g13215,g13188,g13175,g11147,g8238
	,g14521,g14547,g7598,g12644,g12878,g12882,I13805,g10805
	,g11183,g12836,I14765,g13869,g13297,g14231,g13997,g14573
	,g9912,I15042,I13779,g9310,g14741,g14817,I14800,I14482
	,g12870,g11471,g11576,g14333,g12910,g10804,g13870,g14872
	,g12686,g13855,g13384,g12888,g14215,g7201,I14205,g9528
	,I14259,g12860,g12841,g13521,g13300,g13851,I15175,g14793
	,g14754,g12907,g7897,g13886,g10532,g10620,g10509,g10606
	,g10607,I14192,I14346,g10487,g10597,g10572,g10612,g10613
	,g12820,g10571,g14713,g11428,g14772,g12462,g12930,g13120
	,g13140,g13173,g13239,g13255,g13132,g13209,g13142,g13176
	,g13137,g10417,g12026,g12487,I14602,I14650,I14690,g12337
	,I14633,I15831,I16917,g11402,g12845,g12842,g13102,g10816
	,g13501,g10815,g12872,I15342,g14567,g13289,g9908,g14209
	,g14405,g11325,g11498,g14643,g12760,I14611,g11048,I14352
	,g13504,g13295,g14186,g12874,g14914,g11371,g13632,g14432
	,g13663,g13596,g13763,g13625,g8359,g13797,g11367,I15295
	,g11164,g12705,g12972,g11410,g11468,I14708,g12378,g12543
	,I14653,g12598,g13972,g13779,g13676,g14029,g13914,g12818
	,I14579,I14623,g10531,g10503,g10419,g12868,g13217,g13063
	,g11560,g14413,g12640,g11608,g11403,g12137,g12906,g12590
	,g12211,g14503,I15254,g14489,g14520,g14615,g13296,g13939
	,g13910,g12155,I14668,I14687,I14727,I14761,g11032,g11373
	,g14993,g14688,g14691,g14727,g12936,g14434,g14899,g15024
	,g14974,g14776,g12834,g7869,g13871,g13411,g12880,g14416
	,g12937,g9258,g13095,I13872,I14660,g12790,g11404,I14277
	,g12922,g11868,I14630,I14705,I14730,I14647,I14702,I14684
	,I14644,I14671,g11819,g12491,g12819,g10737,g11652,g14601
	,g14062,g14638,g14504,g9825,g14251,g13346,I14248,g12844
	,g14588,g11290,g14613,g12672,g12893,g11234,I14885,g12837
	,g11709,g14515,g14395,g8737,g13301,g13885,g13594,g14364
	,I14749,I14830,g9830,g14537,g14272,g13976,I14899,g14565
	,g12629,g14908,g10887,g14641,I15255,g12861,g13046,g12892
	,g13491,I14663,g11686,g10530,I14589,g10418,g11324,g13378
	,g12929,I16010,g12811,g14535,g14342,g14376,I16898,g7885
	,g12840,g14950,g14984,I14992,g13483,g13141,g14751,g14449
	,g10554,g10475,g13715,g13679,g13621,g13655,g11930,g14275
	,g13637,g13675,g13620,g13593,g11431,g11202,g12895,g12921
	,g14197,g10498,g10812,g8913,g11547,I15800,I14351,g11268
	,g13133,I15043,g12656,g9750,I15129,I15316,g10830,g12975
	,I14993,g12894,I14745,g12914,g12881,g11663,g12614,g11215
	,g14406,g11425,g11615,g13506,g14377,I15176,I16024,g13565
	,g10570,g13626,g10502,g13026,g10474,I14576,g13707,g10776
	,g10685,g14226,I13759,I13762,g12873,I14016,I14069,I14006
	,I16231,g12793,I14305,g10857,g14393,g12911,g12414,g14731
	,g14726,I14854,I15130,g14394,I14610,g14378,g14146,g13945
	,I14290,g14568,g13266,g13248,g13283,g12971,I14714,I15299
	,I14517,g14367,g14339,g13038,I14206,I14170,g13513,I14924
	,g14642,g13524,g13077,g13597,I14766,g13850,g14600,g14574
	,g12342,g14687,g12093,g12511,g12029,g14611,g14505,I15307
	,g14585,I15364,I15335,g14396,g13706,g14538,g14121,g14337
	,I15213,g13436,I14734,g13989,I14855,g14003,g13996,g13971
	,g14089,g14317,g12524,g14821,I15300,g13525,g14360,g14767
	,I14509,g13884,g13025,I16111,g13091,g11185,g13660,g13623
	,g14444,g14447,g10754,g14344,g14911,g14712,g14450,g14831
	,g14033,I15122,g14513,g15042,g14947,g14782,g15033,g14905
	,g15039,g14546,g12933,g14391,g13287,g14433,g11405,g12123
	,g12377,g10775,g13383,g13854,g13542,I14957,g14180,g10476
	,g13495,g13509,g14640,g14362,g14445,g14176,g14516,g14539
	,g13947,g14397,g10590,I15079,I15052,I14789,g14092,g13970
	,g13937,g13712,g13742,g14540,I15123,g14419,g14036,g14001
	,I14735,g14122,g13512,g13796,g13568,g13728,g13820,g14163
	,g12925,g13852,g13202,g13908,g13672,g13883,g13709,g14181
	,g13919,g14637,I15264,g13764,g14832,g14091,I15287,I16721
	,g13666,g14679,g13822,I15937,g14334,I16747,I14230,g14037
	,g14678,g11626,g13990,g13960,g13929,g14154,g14168,g13385
	,I14818,g14064,g13667,g13105,I13852,g14675,g14707,g13600
	,g14697,g14768,g14996,g14732,g12609,g14610,g13324,g13940
	,g14626,g13823,g13143,g13124,g13093,I14229,g13473,g14379
	,g13284,I13851,g13060,g14093,g14708,g14773,g15021,g12667
	,g14548,g14572,g14448,g12954,g13307,g13846,g13260,g13508
	,g10838,g12450,g14761,g14764,g14804,I14518,I15089,g13944
	,g14414,g13736,g14343,g13047,g11492,g11255,g10756,g11225
	,g13665,g14000,g14512,g12924,g13867,g14258,g13518,g14514
	,g14431,g14194,g14027,g14797,g14720,I14427,g14599,g12947
	,g14228,g13294,g11590,g13994,g12920,g14164,g14253,g13946
	,g13246,g13216,g13190,g13342,g13116,g14365,g11890,g13657
	,I14291,g12641,g11432,g13948,g13951,g13977,g14095,g13821
	,g14223,g13247,g12981,g14130,g14110,g13983,g13898,g14133
	,g14015,g14420,I15105,g14090,g14188,g14145,g14278,I16129
	,g13938,g13664,I15080,g14279,g13480,I15214,g13761,g14682
	,g13349,g13281,g14875,g14913,I14925,I15053,g13861,g11144
	,I14790,g14655,g13333,g13762,g13798,g14120,I15365,I15308
	,I14171,g13835,g14366,g13680,g13745,g12932,g14338,g13144
	,g14315,g13782,g12983,g13605,g13416,g13716,g13638,g14336
	,g14591,g14290,g13329,g13394,g13177,g14314,g14398,g12955
	,g13350,g13809,g14454,g13191,g14363,g12857,I17989,I18060
	,I18063,I17956,I17842,I17876,I17916,I18117,I17839,I17754
	,g13017,g13074,g12977,g13027,g13010,g14252,g13041,g13009
	,g14330,g12946,g13101,g14383,g13018,g14276,g12978,g13012
	,g13003,g13055,g12951,g13011,g13075,g12938,g13028,g12918
	,g12976,g11237,I16489,g17134,g13943,g10710,g10851,g10727
	,g10348,g10347,g15819,g14107,g14072,g16610,g15804,g14261
	,g12286,g11761,g11705,g13603,g13574,g11906,g12336,g16672
	,g17119,g11153,g16199,g16535,g15880,g17177,g14320,g13853
	,I17460,I15862,I15194,g15851,g12953,g16705,g11944,g13897
	,g11929,g16593,g16673,g17315,g14522,g14425,g15837,g12136
	,g12490,g15967,g14569,g12538,g16670,g14035,g15815,g12187
	,g13004,g11323,g13223,g13969,g14988,g13156,I16593,g15783
	,g15848,g16841,g16187,g13539,g16516,I16163,g15859,g16871
	,g16424,g15793,g17057,g11559,g15818,g15568,g15030,g17791
	,g15011,g15829,g14247,I17446,g17617,I18421,g13092,g17243
	,g17693,g14873,g16736,g16642,g13005,I16512,g13129,g12979
	,g13545,g16532,g17784,g16596,g11720,I18680,g11845,g12431
	,I18492,g14348,g17777,g14978,g14785,g15045,g14347,I18385
	,g12039,g15669,g16844,g12931,g15808,I17379,g11986,g16730
	,g11931,I14497,g14830,g13778,g12028,g13377,g15823,I15869
	,g16292,I15242,g12100,g13968,I15981,g11189,I18633,g16305
	,g16590,g13282,g13030,g17586,g13139,g12980,g11855,g11820
	,g11872,g11894,g11823,g11920,g11897,g11790,I16120,g11206
	,g13094,g16484,g16614,g15840,g14946,g11842,g10499,g16483
	,g17718,g17585,g17648,g17505,g13044,g17521,g17642,g14924
	,g14882,g17498,g17603,g13013,g16173,g11941,g11917,g11875
	,g11852,g14204,g16926,g16612,g17412,g13325,g13110,g13479
	,g16637,g13415,g13125,g13341,g14309,g15810,g13114,I16596
	,g15705,g13021,g14014,g14422,g16757,g11772,g11706,g16876
	,g16261,g11829,g11900,g15647,g17741,g12436,I15834,g12477
	,g14211,g13833,g16537,g15614,g10488,g13414,g13312,g14034
	,g13305,g14063,g14179,g13458,g13323,g13999,g14032,g13474
	,g14584,g13334,g13975,g14166,g14065,I16468,g14636,g14750
	,g16808,g17138,g12539,g15106,g17213,g15872,g11980,g16758
	,g14912,g13267,g11793,g11878,g11826,g11744,I16733,g13737
	,I16538,g13104,g15912,g16185,g11317,g11136,g11193,g14437
	,g10589,g15995,g15813,I14399,g13907,g16591,g11511,g14216
	,g11966,g17609,g17527,g10363,g15812,g15820,g16518,I15846
	,g13040,g10385,g15727,g16663,I13889,g11294,g17474,I15148
	,g17496,g17600,g14876,g18061,g14794,g17673,g17414,g17518
	,g13290,g11135,g16706,g16608,g16725,g16529,g16658,g17746
	,g17721,g17611,g17651,g13086,I16492,g17416,g17522,g14962
	,g17579,g14845,g17476,g12224,g14496,g13517,g15608,g16731
	,I18417,g15861,g10384,I14369,g13516,I14370,g13942,g14066
	,g16582,g16652,g16522,g16623,g14038,g17681,g17524,g17479
	,g17606,g13824,g13772,I15811,I18449,I16471,g12183,g17153
	,g13189,I15821,g16774,g17144,g16704,I18452,I14400,g13584
	,g13932,g16773,g16630,g16814,g16589,g16692,g14382,g16280
	,g15830,I16676,I16028,g14149,g14205,I15921,g14183,I15954
	,g14169,I15918,g14150,I15932,g14203,g14191,g14184,I15942
	,g14219,g14255,I15987,g12144,g13278,g13061,g13106,g13082
	,g13484,g13036,g13037,I16610,g13505,g13062,g13522,I16663
	,I15727,g13117,I16579,I16660,I16688,g13498,g17726,I15878
	,I16564,g17612,g17589,g15755,g17473,g17390,g16842,g13109
	,g17738,g15479,g14803,g14187,g14297,g17737,g17583,g14700
	,g17756,g17645,g17503,I16289,g16030,I15166,g14598,g11987
	,g13174,g15746,g13974,g17771,g15756,g16311,g15814,I14530
	,g16843,g14088,I16651,I17474,g16581,g17735,g15344,g14664
	,g16583,g14104,g16472,g16509,g14005,g16602,I15872,g16771
	,g17124,g17499,g17477,g17762,g15842,g16515,I15814,I14211
	,g13555,g14136,g13901,g14045,g16743,g17676,I15243,g14581
	,g16634,g14411,g13888,I17416,I15843,g10473,I17883,g14271
	,g15794,g12077,g12858,g12108,g16689,g16655,g16585,g16527
	,g13515,g14528,g14555,g17759,g15562,g13887,g15731,g17137
	,g16645,g16869,I15765,g14238,g17497,g14630,g17389,g17472
	,g17576,g17707,I13906,g11336,g16482,g15750,g16617,g13631
	,g16740,g17092,I15149,g16720,g16523,g16510,g16584,g16605
	,g14321,g17610,g17758,g14744,g17684,g17774,g17528,g17571
	,g16076,I14428,g17194,g15856,g15805,g16531,g15882,g14971
	,g15027,g13118,g14740,g13321,g14387,g13738,g13832,I15195
	,g12370,g14452,g14054,I18536,g17420,g12221,g16635,g15721
	,g17312,g13084,g16759,g14781,g13131,g16702,g13633,g14706
	,g16047,g14838,g14921,g16519,g15821,g14517,g13866,g16282
	,g16639,g16760,g17418,g17682,g16245,g17748,g16804,g13335
	,g17753,g16066,g15992,g16027,g15786,g16190,g13097,g15850
	,g15796,g16176,g15779,g15807,g15591,g14529,g14575,g16805
	,g13622,g13697,g16233,g16866,I15106,g17405,g17321,g16513
	,g13031,g14854,g13319,g17469,g15825,g16811,g15914,g16728
	,g13100,g14987,I15107,g16422,g17810,g17719,g15803,g14696
	,g16802,g16616,g15704,g16090,g16072,g17146,g15792,g15594
	,g13098,g16803,g15749,g16970,I15288,g16512,g16626,g16526
	,g16742,g16606,g16511,g16281,g15841,g12066,g16258,g16296
	,g16669,g13499,g15784,g13808,g12191,g17596,g16288,g14123
	,g13320,g10543,g13299,g14898,g16208,g14570,g15913,g16684
	,g16268,g16243,g13069,g13604,g16473,g16717,g16716,g13876
	,g13530,g11224,g14674,g13076,g17364,g14590,g13928,g16674
	,g17401,g16764,g17493,g13056,g13830,g13108,g13912,g16260
	,g16696,g15732,g17363,g13042,g17655,g15740,g13050,g16734
	,g14519,g16619,g16986,g13529,g13671,g13661,g13698,g13067
	,g16930,g17643,g13882,g14542,g17424,g16506,g17480,g16766
	,I14330,g17123,g13807,g14930,g15002,g17284,g16592,g15628
	,g16761,g17713,g16536,g11962,I14429,I17494,I18587,g17672
	,g17415,g16239,g15875,g17654,g13119,g16870,g14497,g14549
	,g13078,g15585,g16699,g15965,g16867,g13700,g13765,g14399
	,g13462,g14490,g16690,g13032,g17307,g16221,g16737,g14113
	,g14160,g17239,g15883,g16534,g16746,g15809,g12969,g16671
	,g13066,g16653,g17149,g16667,g17601,g13313,g14889,g14965
	,g16022,g13771,g13730,g13799,g16021,g15712,g16965,g13020
	,g13306,g17574,g16211,g11561,g17417,g17710,g17709,g14668
	,g14262,g17769,g14079,g14139,g16313,I17404,g14583,g16882
	,g16290,g16182,g15747,g12939,g17506,g17246,g16259,g13029
	,g11737,g16707,g13564,g17391,g16638,g17500,g17317,g17292
	,g14306,g16896,g15005,g14937,g17504,g17584,g17189,g16052
	,g17309,g13393,g10472,g15739,g16306,g16839,g13083,g11169
	,g16586,g13526,g15754,g17523,g17478,g17582,g17502,g16641
	,g13497,g14291,g15715,g15831,I18579,I17923,g16528,g16588
	,g16607,g16629,g14639,g13437,g16524,g16299,I15289,g16303
	,g16507,g17482,g15655,g17811,g15707,g11923,g14556,g14602
	,g17220,g12285,I18543,g13461,g16611,g16598,g17396,g16321
	,g13249,g13222,g17492,g12592,g13858,g16618,I18495,g13998
	,g17399,g16883,g12999,g14681,g14719,g14654,g13463,g13107
	,g13485,g13065,g16959,I16755,g14714,g14541,g14833,g16885
	,g12482,g16448,g17637,g17529,g17776,g17652,g17588,g17530
	,g17687,I18485,g15700,g16202,g17595,g15910,g13478,g16928
	,g12478,g14608,g12001,g16800,g13221,g14511,g17525,g17225
	,g16075,g16927,g11118,g15968,g17494,g17467,g14977,g14078
	,g15017,g14936,g14888,g14044,g14844,g14119,g17573,g15678
	,g15574,g15710,g16278,g16238,I18625,g16476,g15738,g13277
	,g17198,g17190,g17393,g16517,g17217,g15582,I18529,g15817
	,g16595,g16324,g16430,g16597,g16304,g15822,g14193,g14210
	,g17692,g16613,g14227,g15839,g15508,g15372,g16636,g13500
	,g17786,g16621,g16474,g16729,g17156,g16316,g16275,g17174
	,g17148,g16319,g17287,g15871,g17290,g15881,g15838,g14625
	,g13670,g15170,g17954,g13805,g15870,g16044,g16197,g15578
	,g15570,g15795,g13656,g15699,g15117,g15120,g15123,g15122
	,g15103,g15114,g15112,g15061,g15118,g15069,g15083,g15131
	,g15146,g15149,g15082,g15098,g15057,g15075,g15150,g15156
	,g15107,g15143,g17657,g15065,g15080,g15062,g15138,g15051
	,g15070,g15147,g15089,g15081,g15068,g15113,g15110,g17727
	,g15054,g17694,g15148,g15073,g15119,g15077,g15128,g15050
	,g15137,g15164,g15115,g15097,g15129,g15121,g18655,g15067
	,g15074,g15124,g15049,g15165,g15056,g15066,g15087,g15141
	,g15079,g15100,g15125,g15053,g15071,g15084,g15132,g15126
	,g15130,g17619,g15152,g15099,g15091,g15092,g15096,g15076
	,g17700,g15090,g15160,g15157,g15144,g15078,g15086,g15142
	,g15154,g15134,g15127,g15060,g15166,g15102,g15116,g15111
	,g15139,g15151,g15161,g15064,g15167,g15155,g15093,g15088
	,g15109,g15072,g15104,g15133,g15135,g15095,g15153,g15094
	,g15101,g15058,g15055,g15162,g15145,g15159,g15059,g15158
	,g15140,g15163,g15108,g15168,g15052,g17663,g15105,g15136
	,g15063,I18301,I18214,I18446,I18248,I18574,I18373,I18280
	,I18526,I18344,I18379,I18310,I17653,I18411,I17750,I18674
	,I18259,I17695,I18364,I18479,I17636,I18367,I18443,I18307
	,I18571,I18408,g16580,g16643,g16963,g16708,g16676,g16644
	,g16738,g16873,g16872,g16767,I17008,I17118,I18168,I18177
	,I18270,I18125,I17763,g17471,g16609,g16631,g17242,g17216
	,g16750,g17411,g16530,g16320,g16726,g17366,g16727,g17301
	,g16695,g16661,g16632,g17470,I18469,I17125,I17198,I18842
	,I17111,I18265,I18143,I18131,I17159,I18120,I17228,I18829
	,I18382,I18313,g17157,I17639,I18078,g17794,I18482,g17489
	,g17465,g17410,I17136,I18865,I17723,I18154,I18104,I18252
	,I18165,I17675,I17401,I17488,I17471,I18083,I17658,I17420
	,I17661,I18849,I17590,I17355,I17098,I17374,I17976,I18028
	,I18048,I18285,I17442,I18003,I18006,I18839,I18852,I18810
	,I18350,I17173,I17679,I17425,I17436,I18101,I17699,I17491
	,I17507,I17154,I17276,I18180,I17249,I18221,I18320,g17512
	,g17491,g17466,I17188,I18832,I18434,I17108,I18875,I18868
	,I17704,I18089,I18151,I18135,I18238,I17101,I17104,I18855
	,I18398,I18822,I17181,I18872,I17392,I18071,I18009,I17456
	,I18031,I18323,I18051,I18034,I17121,I18858,I17128,I18518
	,I17140,I17207,g15858,g16868,g17087,g17147,g17121,g17789
	,g16163,I17447,I17884,I17475,I17380,g15613,g12351,g19209
	,g17736,g12301,g15735,g20172,g20163,g12970,g10544,g16958
	,g17085,g16968,g17733,g13138,g17605,g16023,g16815,g15674
	,g17783,g19356,g17755,I16724,I16698,g19965,I16855,g13279
	,g16732,g15969,g21188,g16694,I20467,g12423,g16688,g16654
	,g16812,g16124,g16158,g16186,I14213,g13251,g20186,g17679
	,g14185,g14221,g16854,g19853,g13304,g16651,g16622,g19611
	,g13057,g14207,g14233,g16024,I17476,g17511,g14536,g15785
	,I20486,I14532,I14531,g15672,g16204,g16668,g17768,I15168
	,g15978,I16629,I15167,g17175,g16183,g17514,g16956,g14031
	,g17086,g17014,g17772,g17135,g17814,g17670,g14316,g14412
	,g13311,g14571,g14543,g14423,g13096,g14544,g14453,g13514
	,g13460,g13431,g13409,g13477,g13410,g13583,g14563,g16200
	,g16853,g16159,g16172,g11389,g13258,g17785,I16775,g14308
	,g15936,g13256,g13211,I18762,I18785,I17542,I18713,g13250
	,g16685,g16423,g17264,g20131,g11350,g15693,g15902,g21430
	,g19576,I18682,g17641,g17602,g14332,g16264,g17599,g17308
	,g10521,I19802,g16845,I15494,g13280,g16846,g15713,I16590
	,g20854,g15725,g16128,g19369,g15507,g16026,g14424,g14753
	,I18635,g19793,g14384,g14616,g12940,g12997,g13016,g12968
	,g16207,g18088,I18879,g16579,I17744,g16222,g20237,g16210
	,g15863,I18620,I18765,I17741,I17552,I18819,I18740,I18568
	,I17585,I18671,I17529,I17606,I17575,I18782,I18716,I18803
	,I17692,g17464,g14307,I16515,g13271,g21510,g13024,g12998
	,g19533,g14443,g15852,g15903,g15876,g17616,g15811,g15799
	,g13007,g13015,g13033,g13045,g20070,g15745,g17677,g17392
	,g14206,I15572,g13793,g12967,g13023,g13034,g12996,g13022
	,g13014,g12995,g13008,g16479,g13510,g19522,g19427,g13303
	,I14499,g16807,I16544,I16626,g16929,g21556,I16679,g17720
	,g17745,g17136,g17122,g17815,g17154,g17569,I16455,I17461
	,g17490,g16215,g16226,g14358,I18370,g20645,I17448,g20870
	,g17763,g17507,g13857,g16227,g16237,g20085,g14442,g16325
	,g16712,g16289,g16680,g16310,g16768,g16739,g15873,I16541
	,g17180,g16198,g13298,g13064,g16721,g16475,I16969,g14331
	,I16160,g16098,g15847,I17324,I17733,I17302,I17772,I17801
	,I17873,I17314,I17834,g15633,g15836,g16177,g16097,g19530
	,g19350,g15701,g15874,g13476,g13496,g13130,g13554,g15653
	,g16161,I18538,g16666,g21333,I17462,g15589,g14256,g16203
	,g16733,g14257,g14220,g16125,I18487,g16687,g15654,g17488
	,g13252,g15718,g17515,g15757,g16220,g16178,g15857,g19614
	,g16765,g19932,g16599,g14295,g16025,g15724,g16193,g19265
	,g21302,g15966,g15717,g19778,g13543,g21253,g19336,I17495
	,I17924,I17405,g14296,I18681,g20187,g19587,g15567,I17381
	,g15673,g13079,I14498,g15864,g15833,g14645,g17809,g15695
	,g15723,g19873,g16485,g16751,g15572,I18634,g13459,g13475
	,g13528,g13115,g17510,g15651,g16184,g15935,g17598,g16806
	,g16701,g19597,g20751,g14222,g16801,g21361,g20871,g15726
	,g16810,g17365,g15706,g17752,g16191,g15937,g17770,g20108
	,g20093,g19605,g17820,g20173,g15853,g15907,g16122,g17297
	,g16231,g17872,g13019,g19344,g18994,g12471,g17792,I18589
	,g16206,g16235,g16214,g17056,g16195,g16223,g16180,g16127
	,g16162,g16099,I18233,g16646,I18581,I18580,g19501,g16201
	,g16966,g16770,g19911,g21389,g21190,I18148,g15849,g20875
	,g20838,g17513,g17717,g17481,g16840,g19467,g16219,g16625
	,I21162,g16633,g17846,g19632,g13413,g16427,g16224,I17406
	,g15679,g16514,g16724,g19274,g16735,g17120,g17754,g17013
	,g16969,g16232,g17734,g17578,g19557,g20202,g16749,g19488
	,g19619,g15709,g16741,g17597,g17419,g17680,g19595,I14332
	,g20272,g16691,g16747,g20217,g21413,g21378,g19518,g21298
	,g19506,g13242,g13264,I18588,I17496,g11419,g16212,g21460
	,g16700,g17644,g17714,I14331,g19475,g17765,g15590,g16287
	,g19275,I19762,g16884,g21285,g16192,g16179,g16171,g16096
	,g16769,g16123,g20276,g19407,g15632,g19857,g19879,I14212
	,g21296,g15753,g17640,g19363,g19362,g19428,g19604,g12239
	,g17708,g17775,g19364,g20241,g19207,I17885,g20887,g17790
	,g17686,g19071,g17268,g19355,g19738,g19408,g20765,g17575
	,g17638,g21347,g19374,g20734,I18537,g16809,g17683,g17742
	,g20212,g21011,g15703,g15722,g17635,g17788,g17757,g16520
	,g16657,g15729,g17716,g15743,g16813,g21140,g15736,g17744
	,g17572,g16875,g17468,g15797,g17647,g19525,g21163,g16723
	,g20739,g15911,g16488,g16538,g17636,g17671,g21024,g17816
	,g17723,g15728,g19359,g17773,g17594,g15612,g17495,g16242
	,g16762,g17145,g16209,g16703,g17570,g15719,g20675,g15652
	,g16772,g16160,g15884,g16925,g19751,g19791,g15860,g15702
	,g20717,g16126,g15720,g20733,g15694,g15611,g16763,g19903
	,g20979,g19916,g15631,g19874,g19887,g21332,g15581,g15744
	,g15716,g21012,g15711,g20676,g15708,g20644,g19795,g19875
	,g21250,g21277,g15962,g15877,g15867,g15844,g20559,I17925
	,g20682,g15782,g19856,g15730,g21206,g17133,I18531,g16855
	,g21124,g17625,g20035,I18486,g20011,g18935,I18627,g21306
	,g20619,g19146,I18626,g19981,g20995,I18530,g15680,g15563
	,g17587,g15483,g17952,g15426,g16826,g16861,g17384,g16821
	,g16077,g16795,g16877,g15915,g18062,g15615,g17818,g17475
	,g17929,g15277,g15224,g17200,g16987,g17059,g16923,g16508
	,g18008,g18065,g15345,g17501,g17844,g15634,g17367,g17183
	,g15733,g17128,g15758,g15573,g16164,g16136,g16489,g16931
	,g16031,g16000,g16449,g15595,g17413,g17812,g17926,g17847
	,g16782,g16777,g16053,g17302,g16856,g16816,g16752,g15885
	,g15171,g15862,g16249,g17873,g16349,g15979,g16326,g16897
	,g16100,g16129,g15938,g16431,g17093,g17226,g16954,g17062
	,g16525,g17955,g15509,g17533,g16886,g16309,g17328,g17433
	,g17821,g15714,g16964,g15579,g16971,g17015,g17249,g15348
	,g17870,g15656,g15480,g17526,g16587,g16967,g17271,g17125
	,g17096,g15373,g15085,I18900,I18903,I18909,I18897,I18888
	,I18891,I18894,I18906,I18885,I18882,g17485,g17614,g17326
	,g17508,g17428,g16308,g17532,g17427,g16487,g17247,g17691
	,g16578,g17486,g16323,g17327,g17432,g17409,g17591,g17296
	,g17430,g17615,g17224,g17509,g17178,g17324,g21652,g21653
	,I20929,I19012,I19235,g21655,I20891,g21656,g21654,I20882
	,I19348,I19487,I19238,I18912,g21658,g21660,I20793,g21659
	,I20840,I20830,g21657,I19345,I19484,g13856,I17094,g15048
	,g19393,g19788,g19691,g19461,g19145,g16662,g13241,g13580
	,g13573,g19589,g19546,g19483,g19513,g16093,I17747,g18910
	,g18933,g19735,g14385,g16279,g20783,g19717,g19736,g20181
	,g22709,g21272,g19948,g17690,g17724,g17613,g17766,g17747
	,g17780,g21251,I17148,g19637,g19660,g13918,g19442,g19588
	,g20094,I18262,g13240,g20188,g16069,g23392,g23391,g17429
	,g20784,g17140,g17176,I17114,g21294,g17699,g14277,g17192
	,g14564,g19564,g19578,g19441,g15904,g14509,g13058,g14386
	,g11545,g20162,g21405,I17780,g19693,g19716,g20171,g20215
	,I17609,g17193,g17662,g13551,g13210,g15832,g16181,g13544
	,g19555,g21403,g19063,g21557,g20169,I18224,g18951,g18981
	,g20107,g12952,g21288,g20375,g20092,g18879,g19510,g19549
	,g19455,g19495,g19267,g19886,g21388,g20160,g19337,g18906
	,I18523,g21377,I20488,g19907,g21354,I17650,g14359,g20165
	,g21301,I18861,g20081,g21331,g16540,g20033,g18091,I19917
	,I17131,g21344,g22983,g20148,g23626,g19450,g14441,g20065
	,g20078,I17671,g12875,g19264,I20468,g19609,g19069,g23079
	,I18376,g21359,g19571,g20199,g17781,g20051,g13877,g21393
	,I17612,g15571,g20063,g21353,I18341,g14676,I17633,g13902
	,I18205,I17808,I17143,g19746,I18476,g12332,g14510,g21360
	,g20007,g14739,g20977,g11591,g20095,I17166,g16119,I17783
	,g20135,g13257,g23292,I17615,g11154,g14745,g19913,g21385
	,g21283,I20469,g20039,I17668,g19474,g14790,g16681,g20203
	,g14582,g14609,g21345,g14695,g17712,g17740,g14771,g19502
	,g21417,g21330,g20055,g20112,I18788,g14730,g20068,g14669
	,g14701,g19962,g19466,g19752,g17150,g17182,g21287,g16719
	,g19139,g19333,g19462,g20082,g17593,g17199,g22859,g23412
	,g23411,g21357,g21416,g15800,g17191,g22304,g20170,g20111
	,g23229,g23151,g13958,g17761,g21394,g20192,g14820,g23055
	,g22870,g22718,g23285,g23132,g22152,g23733,g21363,g14631
	,g13993,g16776,g14780,g19692,g19681,g22760,g22759,g16745
	,g21334,g20077,g20034,g18950,g18993,g18982,g20905,g20193
	,g13043,g21187,g17779,g18974,g19914,g17151,g17091,g21289
	,g13967,I20487,g19061,g19740,g17139,g17152,g21186,g19575
	,g22226,g19358,g21339,g20151,g19266,g20000,g16234,g17817
	,g16539,g16194,g16205,g16213,g21307,g18893,g18909,g19601
	,g19585,g21433,g11292,I20460,g13933,g16155,g17624,g15580
	,g22406,g19997,g19880,g23666,g19354,g22340,g19516,g19521
	,g19767,g13927,g15789,g17179,g23978,g22534,g23659,g20109
	,g13896,g18943,g19535,g17793,g16244,g16283,g17767,g16486
	,g17725,g17653,g19680,g14829,g19536,g15959,I20499,g19335
	,g19449,g19500,g21451,g20218,g19206,g22762,g16893,g22869
	,g23402,g23931,g23645,g17058,g23182,g23051,g20196,g19756
	,g17618,g17181,g16713,g14871,g19487,g20540,g17197,g14786
	,g20388,g20531,g20782,g22871,g19384,g23574,g22680,I20035
	,g19953,g19372,g23424,g23423,g23971,g23714,g22858,g23425
	,g22449,g23711,g22993,g21605,g19524,g20572,g20550,g17568
	,g16957,g19486,g16521,g22217,g23108,g22492,g16196,I22024
	,g16640,g15816,g16675,g16615,g16594,g15806,g16533,g15824
	,g20248,g21062,g19684,g23286,g15843,g18992,g23560,g23678
	,g23309,g17656,g22191,g19784,g23909,g22846,g21348,g21303
	,g23381,g23380,g22172,g17592,g19062,g22753,g23024,g19140
	,g19768,g23756,g22311,g23900,g23208,g18987,g19661,g21284
	,g19749,g19572,g19904,g19593,g19949,g23972,g19855,g20174
	,g17675,g19999,g19715,g19594,g22161,g23729,g19906,g19951
	,g20027,g23890,g19655,g19545,g21365,g23052,g23932,g15650
	,g23602,g23590,g23889,g23563,I23099,g22845,g23382,g22309
	,g22707,g20269,g20328,g20595,g20643,I22769,I22725,g22843
	,g22842,g23103,g22717,g22716,g23726,g18934,g23623,g23401
	,g23400,g14663,g23699,g23681,g23413,g23948,g22896,g22225
	,g23917,g23063,g22654,g23854,g23139,g14686,g23067,g23811
	,g23801,g21351,g23586,g20134,g20185,g22306,g23405,g22669
	,g23779,g23342,g21402,g23112,g22897,g23082,g22761,g23308
	,g22308,g19556,g23630,g22857,g23908,g23605,g23393,g22919
	,g23341,g23127,g22844,g23695,g23949,g21066,g19674,g23642
	,g19656,g23124,g22720,g18890,g18949,g23105,g21382,g22160
	,g21276,g21067,g23692,g23167,g23662,g23135,g18709,g18374
	,g18282,g18343,g18420,g18671,g18656,g19890,g18602,g18305
	,g18774,g18588,g18727,g18756,g18749,g18660,g18494,g18397
	,g18134,g18161,g18641,g18233,g18598,g18505,g18663,g18409
	,g18354,g18676,g18686,g18601,g18315,g18745,g18392,g18520
	,g18171,g18534,g18637,g18604,g18567,g18201,g18616,g18743
	,g18341,g18276,g18603,g18458,g18581,g18783,g18483,g18439
	,g18712,g18269,g18789,g18527,g18106,g18215,g18307,g18633
	,g18698,g18410,g18779,g18612,g19919,g18605,g18569,g18659
	,g18406,g18274,g18230,g18582,g18540,g18757,g20841,g18752
	,g18583,g18333,g18816,g18338,g18472,g18235,g18495,g18524
	,g18335,g18417,g18644,g20014,g18344,g18482,g18138,g18775
	,g18157,g18164,g18454,g18593,g18362,g18212,g18202,g18455
	,g18245,g19402,g18419,g18145,g18462,g18425,g18280,g18340
	,g18543,g18386,g18763,g18631,g18748,g18728,g18767,g21143
	,g18795,g18375,g18185,g18737,g21127,g18786,g18643,g18311
	,g18693,g18708,g18304,g18808,g18391,g18571,g18329,g18390
	,g18563,g18739,g18675,g18370,g18487,g18358,g18741,g18369
	,g20773,g24141,g18773,g18303,g19422,g18691,g18817,g18278
	,g18584,g18302,g18131,g18236,g18500,g18433,g18785,g18347
	,g18211,g18427,g18617,g18228,g18300,g19338,g18824,g18411
	,g18327,g18165,g18592,g20720,g18744,g18268,g18489,g18361
	,g18558,g18266,g18121,g18721,g18553,g18253,g18559,g18506
	,g18424,g18238,g18404,g18275,g18434,g18146,g18324,g18415
	,g18668,g18516,g18535,g20982,g18764,g18365,g18522,g18403
	,g18332,g18760,g18325,g18378,g18259,g18258,g18810,g18342
	,g18104,g18360,g18441,g18436,g18234,g18112,g18163,g18160
	,g18277,g18367,g18541,g18576,g18471,g18547,g18449,g18428
	,g18717,g18484,g20781,g24144,g18435,g18478,g18822,g20857
	,g18761,g18536,g18126,g18765,g18267,g18459,g18376,g20705
	,g18285,g18753,g18806,g18799,g18653,g18317,g18408,g18646
	,g18568,g18431,g18298,g18490,g18176,g21209,g18812,g18718
	,g18349,g18218,g18359,g18371,g18107,g18372,g18150,g18412
	,g18210,g18530,g18513,g18479,g18623,g18262,g18184,g18826
	,g18538,g18270,g18544,g18456,g18246,g18713,g18678,g18523
	,g18273,g18542,g18477,g18466,g18742,g18400,g18680,g18232
	,g18102,g18768,g18734,g18265,g18389,g18443,g18159,g18260
	,g18162,g18590,g18797,g18183,g18706,g18531,g18720,g18504
	,g18447,g18414,g18480,g18488,g18366,g18578,g18205,g18174
	,g18762,g18147,g18193,g18263,g18192,g18208,g18158,g18554
	,g18321,g18142,g18401,g18206,g18642,g18724,g18674,g18595
	,g18689,g18736,g18758,g18533,g18153,g18529,g18444,g18615
	,g18609,g18701,g18445,g18792,g18387,g18256,g18751,g18501
	,g18295,g18515,g18492,g18364,g18152,g18546,g18399,g18658
	,g18465,g18216,g18463,g18328,g18499,g18682,g18254,g18182
	,g18220,g18127,g18719,g18572,g19968,g18622,g18385,g18297
	,g18384,g18136,g18448,g18497,g18725,g18549,g18379,g18248
	,g18574,g18813,g18306,g18151,g18575,g18688,g18532,g19984
	,g18636,g18286,g18320,g18591,g18791,g18141,g18502,g18491
	,g18723,g18293,g18197,g18667,g18299,g21256,g18815,g18818
	,g18526,g18191,g18155,g18577,g18377,g18521,g18684,g18240
	,g18608,g18606,g18811,g18638,g19935,g18619,g18733,g18825
	,g18519,g18460,g18422,g20998,g18778,g18692,g18679,g18654
	,g18405,g18196,g18771,g18630,g18187,g18669,g18430,g18645
	,g18166,g18115,g18759,g18661,g18363,g18699,g18330,g18819
	,g18398,g18467,g18685,g18780,g18125,g18452,g18509,g18128
	,g18382,g18284,g18528,g18700,g18566,g18662,g18251,g18690
	,g18113,g18772,g18139,g18292,g18508,g18137,g18129,g18620
	,g18334,g20915,g24139,g18510,g18237,g18279,g18555,g18730
	,g18170,g18468,g18429,g18517,g18350,g18322,g18241,g18512
	,g18143,g18626,g18446,g18351,g18635,g18110,g18790,g18103
	,g18613,g18625,g18556,g18116,g18589,g18199,g18189,g18395
	,g18252,g18119,g18657,g18156,g18514,g18373,g18696,g18353
	,g18475,g20922,g18611,g18801,g18135,g18496,g18507,g18225
	,g18314,g18402,g18551,g18453,g18407,g18777,g18432,g18687
	,g18461,g18747,g18383,g18264,g18213,g18704,g18539,g18561
	,g18132,g18336,g18421,g18470,g18493,g18639,g18738,g18357
	,g18814,g18261,g18118,g18537,g18120,g18481,g18290,g18648
	,g18221,g18242,g19268,g18579,g18705,g18310,g18464,g18289
	,g18511,g18796,g18597,g18308,g18423,g18766,g18457,g18316
	,g18437,g18313,g18223,g18570,g18249,g18781,g18665,g18124
	,g18607,g18130,g18707,g18672,g18649,g18250,g18326,g18621
	,g18200,g18820,g18677,g18651,g18178,g18108,g18272,g18416
	,g18545,g18281,g18729,g18585,g18769,g18355,g18203,g18552
	,g18440,g18793,g18473,g18231,g18255,g18331,g18111,g18629
	,g18803,g21193,g18650,g18548,g18219,g18754,g18204,g18190
	,g18226,g18722,g18800,g18640,g18476,g18368,g18681,g18485
	,g18418,g18227,g18173,g18396,g18697,g18123,g18807,g18784
	,g18318,g18627,g18586,g18109,g18168,g18105,g18565,g18550
	,g18442,g18726,g18732,g18614,g18573,g18610,g18740,g18735
	,g18469,g18244,g18782,g18337,g18294,g18474,g18243,g18702
	,g18426,g18301,g18710,g18823,g18587,g18628,g18271,g18186
	,g18288,g18770,g18525,g18673,g18287,g18695,g18175,g18393
	,g18346,g18312,g18794,g18291,g18296,g18323,g18144,g18694
	,g18715,g18179,g18596,g18352,g18207,g18486,g18746,g18172
	,g18133,g18755,g18809,g18239,g18802,g18167,g18247,g18750
	,g18224,g18714,g18214,g18560,g18594,g18600,g18154,g18664
	,g18194,g18169,g18394,g18683,g18380,g18716,g18229,g18198
	,g18599,g18209,g18257,g18149,g18148,g18634,g18787,g18731
	,g18413,g18804,g18180,g18222,g18564,g18309,g18283,g18451
	,g18821,g18666,g18703,g18503,g18618,g18805,g18798,g18181
	,g18122,g18518,g21061,g18670,g18388,g18345,g18632,g18438
	,g18339,g18319,g18624,g18177,g18711,g18652,g18217,g18195
	,g18788,g18188,g18356,g18348,g18580,g18776,g18117,g18114
	,g18140,g18498,g18647,g18450,g18381,g18557,g19638,g19417
	,g19376,g19757,g19773,g21222,g19620,g19345,g19626,g19662
	,g19379,g21370,g18984,g20204,g20097,g21156,g20277,g18954
	,g19389,g20242,g21225,g21160,g19330,g19606,g21308,g18093
	,I19384,g18876,g20503,g21408,g21274,g21422,g20609,g20664
	,g21179,g20914,g20665,g21054,g20704,g20383,g20444,g20545
	,g18887,g21052,g20634,g20564,g20663,g21454,g20913,g21053
	,g20703,g20587,g20502,g19800,g19677,g19861,g20238,g19771
	,g19732,g19712,g19687,g19742,g19787,g19743,g20025,g19996
	,g20533,g20026,g19878,g20040,I20937,I20584,I21210,g20555
	,g21204,g21205,g21252,g20737,g18880,g21155,I19796,g20625
	,g20514,g20435,g20538,g20554,g20680,g20650,g20498,g20600
	,g21461,g19885,g20903,g20004,g20656,g20087,g20579,g20179
	,g19747,g20247,g19695,g20207,g19776,g19629,g19777,g19718
	,g19649,g19760,g19682,g19789,g19761,g19852,g19748,g20229
	,g19696,g19737,g20320,g19872,g19790,g20190,g19698,g20167
	,g20158,g19650,g20178,I21006,I20913,I21115,g20191,g20541
	,g21346,g21355,g20379,g20209,g21418,g20523,g20265,g20321
	,g20231,g20103,g20766,g20005,g20036,g20657,g20697,g20627
	,g20104,g20090,g21049,g20105,g19960,g20904,g20601,g20066
	,g20067,g20147,g20106,g20560,g20053,g20037,g20079,g20080
	,g20129,g20091,g20006,g20130,g19961,g20580,g19912,g20038
	,g20054,I20529,g20157,g20166,g19697,g20102,g20088,g20089
	,g20146,g20052,g20064,g20101,g20144,g20159,g20696,g20145
	,g20128,g21048,g20208,g21295,g20168,g20180,g20671,g21182
	,g18889,g21249,g20591,g21183,g20507,g21286,g20712,g21456
	,g21060,g21059,g20529,g20448,g18897,g20779,g20710,g20780
	,g21184,g20711,g20641,g20530,g21466,g20615,g20568,g21425
	,g21380,g20562,g21396,g20629,g20701,g20324,g20770,g18828
	,g20605,g20585,g21178,g20501,g20630,g20267,g20525,g20380
	,g21406,g20768,g20769,g21608,g20702,g20381,g20606,g20607
	,g20543,g20909,I20562,g19676,g19659,g19754,g19770,g19799
	,g19686,g20213,g19730,g19786,g19711,I20895,g19979,g19860
	,g19980,g19947,g20010,g20510,g19731,g19409,g19763,g19395
	,g19477,g19386,g19387,g19779,g19396,g19468,g19451,g18883
	,g18874,g21604,g18944,g19558,g18884,g18975,g19537,g19539
	,g19577,g19559,g19523,g18946,g19273,g19538,g18976,g18977
	,g18945,g18929,g18908,g19670,g19612,g19719,g20194,g19652
	,g19653,g19630,g20182,g19765,g20110,g20210,g19762,g19469
	,g19385,g19394,g19434,g19421,g19963,g19476,g19368,g19452
	,g19750,g18885,g19067,g18907,g18988,g19542,g19437,g19493
	,g19586,g19569,g19543,g19618,g19480,g19526,g19503,g19527
	,g19481,g19472,g19491,g20009,g19473,g19414,g19570,g19454
	,g20057,g19494,g19915,g19617,g19544,g19657,g19602,g19528
	,g19529,g19504,g19603,g19505,g19482,g19634,g19492,g19635
	,g21050,g21379,g20659,g20700,g20698,g20699,g20767,g20604
	,g21607,g20500,g21362,g20584,g20441,g20524,g20266,g20561
	,g20322,g20323,g21395,g20603,g20582,g20233,g20583,g20542
	,g21560,g20660,g19431,g19360,g19438,g19365,I20216,g20526
	,g20910,g20661,g20632,g20911,g21051,g21397,g20633,g20563
	,g20325,g18829,g20771,g20608,g20382,g18875,g20544,g20631
	,g21247,g21421,g20662,g21407,g20912,g20442,g20586,g20772
	,g20443,g19905,g19416,g19366,g19950,g19744,g19439,g19865
	,g19432,g19678,g19498,g19531,g19713,g19733,g19552,g20551
	,g20059,g18916,g18938,g18904,g18891,g18952,g19517,g19688
	,g20058,g20096,g19679,g19499,g20153,g19553,g20597,g20240
	,g20535,g20494,g20432,g20552,g21400,g20574,g20274,g20372
	,g20495,I19756,I21181,g20978,g20732,g20852,g20622,g20853
	,g21561,g19373,g19479,g19410,g19443,g19766,g20008,g19435
	,g19489,g19471,g19780,g19397,g19565,g18978,g18894,g19579
	,g18895,g19478,g18886,g18989,g19470,g18827,g18931,g18896
	,g19144,g19068,g20211,g19654,g19739,g19633,g20195,g19683
	,g20132,g20232,g19783,g19672,g19673,g19781,g19411,g19490
	,g19794,g19398,g19399,g19429,g19412,g18979,g18980,g18990
	,g18947,g18991,g19541,g19566,g18932,g19343,g19600,g19580
	,g19567,I21067,g21428,g21412,g18903,g19415,g19352,g21349
	,g21305,g21467,g21458,g21337,g20273,g20239,I20690,g19772
	,g20534,g19208,g19351,g21457,g21427,g19276,g21304,g21383
	,g21336,g18832,g20679,g21138,g21139,g21189,g21010,I19786
	,I21199,g20537,g20624,g20497,g20649,g20434,g20576,g21431
	,g20374,g20599,g20513,g20536,g20706,g20384,g20707,g20527
	,g20546,g20385,g20776,g20612,g21381,g21409,g20636,g21180
	,g20588,g20610,g18830,g20774,g20611,g20775,g20504,g21398
	,g21609,g20326,g20635,g20565,g20268,g20916,I20542,I20846
	,g19710,g20197,g19685,g19741,g19658,g19785,g19636,g19675
	,g19709,g19753,g19769,g19964,g19930,g19931,g19902,g19798
	,g20452,g20917,g18877,g20547,g21248,g20446,g20777,g20613
	,g21423,g20566,g21410,g20637,g20589,g21055,g20918,g20919
	,g20528,g20445,g18831,g20386,g20778,g21399,g20327,g20638
	,g20639,g20666,g20667,g20923,g20450,g20714,g20715,g20451
	,g20389,g20235,g20329,g20674,g20594,g20570,g20642,g20616
	,g20617,g20270,g20713,g21426,g20571,g20532,g20549,g20716
	,g20449,g20672,g20592,g20508,g20509,g20673,g21185,g20593
	,g20569,g20618,g21068,g21069,g20496,g20623,g20598,g20433
	,g21414,g20553,g20575,g20275,g20373,g20511,I21189,I19772
	,g20648,g21123,g20994,g20869,g21610,g20993,g20512,g19952
	,g19370,g19440,g19755,g19445,g19433,g19998,g19881,g19573
	,g19745,g19689,g19519,g18917,g18939,g18905,g18983,g18953
	,g19714,g19532,g20573,g20072,g19734,g19554,g20071,g19520
	,g20113,g20164,g19690,g19574,g21057,g20590,g18888,g20447
	,g20506,g20920,g21275,g20921,g20567,g21411,g20668,g20669
	,g21181,g21058,g20708,g20709,g18878,g20548,g20387,g20505
	,g20640,g20614,g21455,g21424,g20670,g21056,I19813,g20738
	,g20515,g20539,g20577,g21511,g20499,g20626,g20681,g20651
	,g20556,I19661,g20578,g21279,g21268,g20874,g18892,g21221
	,g21267,g20152,g20084,g23770,g22640,g17581,g24140,g17782
	,g21895,g21894,g16628,g23217,g21401,g17705,g17669,g23436
	,g23885,g17650,I17919,I17626,I18304,g16428,g20201,g15781
	,g21415,g16286,g24280,g21892,g17668,g22644,g23920,g16601
	,g23298,g23348,g15737,g20234,g19436,g23318,g15588,g20216
	,g21897,g21900,g23957,g23346,g22158,I17557,g17531,g23358
	,g15566,g16620,g17155,g16307,g20581,I18245,g17408,g24142
	,g21464,g16285,g17634,I19778,g17431,g21558,g21404,g22662
	,I21722,g16429,I18160,g24999,g23324,g19560,g23856,g16246
	,g19631,g20184,g15506,g19446,I21222,g21690,g20060,I21258
	,g19908,g21662,g19866,g19957,g21666,g21694,g21670,I21230
	,I21242,g19882,I21250,g21682,I21226,g19954,I21246,g20046
	,g21674,g19869,I21234,g20073,g21686,g21678,I21238,I21254
	,g21893,g17953,g21420,I18414,g16322,g21901,g17590,g22359
	,g22407,g22529,g22496,g22457,g22369,g23234,g19540,I17395
	,g17188,g22384,g22649,g22547,g16272,g16284,g24143,g16600
	,g22331,g21899,I17879,g15748,I18114,g23194,I17569,I18138
	,g23919,g15371,I21047,g23319,g17248,g15569,I19775,I21058
	,I21074,I20355,I20388,I20369,g21891,I18191,g23345,g22625
	,g16577,g22497,g22408,g22527,g22544,g22679,g23296,g15169
	,I18086,g23251,g23204,g23042,g20522,g24787,I21042,I19831
	,I21013,I19843,I19851,I19863,I21029,I19857,g22645,g19596
	,g24378,g16312,g22863,g22719,g24482,g16236,g23276,g19388
	,g16604,g19651,g20390,g19430,g23261,g24649,g19610,g22653
	,g24014,g22312,g19383,I20461,g24416,g25448,g23297,g23884
	,g24603,g19444,g23836,g25237,g22216,g23047,g20628,g23855
	,g23197,g24011,g16291,g19401,g23822,g22588,g22530,g24720
	,g24640,g16225,g24008,g22342,g22417,g22472,g24796,g22209
	,g20183,g19400,g23720,g15741,g22901,g22432,g22498,g19592
	,g23153,g23171,g23087,g24785,g25160,g21453,g21606,g21465
	,I20910,g22193,g23129,g23383,g24758,g22665,g23716,g24545
	,g24607,g15734,g22708,I22918,g22298,g24687,g22751,g20230
	,g24766,g21452,g21419,g17520,g24820,g24953,g25366,I19704
	,I19734,I20569,I19759,I20495,I20447,I19789,g22641,g23615
	,g22685,g23850,g25273,g18930,g23374,g25285,g24580,g24731
	,g25109,g25001,g25092,g25016,g22664,g19453,I16778,g23209
	,g22591,I20412,I20399,I20385,I20609,I19799,I20433,g22860
	,g15752,g15787,I23149,g20214,g20149,g19413,g23795,g23331
	,g20658,g25047,g25153,g25036,g25133,g24809,g21432,g15742
	,g15780,g17608,g22318,g15751,g18948,g22684,g22832,g20198
	,g25034,g24730,g24387,g19581,g20602,g24430,g25216,g22307
	,g22208,g25072,g24987,g25000,g25090,g23193,g23183,g22219
	,g24903,g23062,g24557,g24790,g24659,g22299,g24604,g24683
	,g24587,g24667,g21462,g19613,g24590,g24776,g16660,g17732
	,g24398,g19671,g22937,g24628,g22639,g24484,g23007,g24922
	,g24421,g24795,g22648,g24390,g17706,g23275,g24565,g15798
	,g24528,g25229,g22634,g24411,g24713,g24985,g23262,I20462
	,g21513,g24401,g24443,g19568,g22636,g24475,g24665,g24586
	,g24579,g24655,g23009,g24670,g24582,g17689,g23871,g24930
	,g21384,g25172,g24501,g24605,g24626,g24711,g24685,g25255
	,g20083,g20076,g24437,g23104,g24585,g25035,g25131,g25111
	,g25017,g25186,g24415,g23750,g23050,g25233,g24608,g24701
	,g22218,g25293,g24940,g25037,g15788,g23578,g23620,g24395
	,g24403,g23954,g24986,g25070,g25055,g24971,g19534,g25202
	,g23255,g25174,g25046,g25327,g23317,g22325,g22142,g24432
	,g25203,g23835,g25239,g22991,g22659,g23782,g22939,g19070
	,g25334,g22660,g23023,g22538,g25188,g24789,g22652,g24778
	,g23472,g23130,g23512,g23192,g23530,g23614,g23654,g23550
	,g23496,g23573,g24392,g24436,g24569,g25144,g25189,g24488
	,g24625,g24450,g24771,g25015,g23883,g24671,g24588,g24913
	,g24629,g24581,g22190,g24686,g24814,g24572,g23686,g24589
	,g24606,g25268,g24639,g24409,g24714,g24556,g24757,g24422
	,g24751,g24464,g23918,g24410,g24399,g24465,g24400,g24423
	,g24393,g24550,g23955,g24804,g24842,g24793,g24451,g25200
	,g24495,g24402,g24427,g25218,g25175,g24779,g23763,g18833
	,g19277,g19074,g21514,g22310,g20785,g20330,g21562,g19147
	,g20596,g21335,g21468,g18997,g19801,g20924,g20391,g23280
	,g20283,g23220,g21387,g21037,g21273,g19210,g21611,g20453
	,g21070,g18562,I22729,I22485,I22665,I21792,I21802,I21757
	,g23223,g23211,I21815,g23844,g23789,I21776,g23239,g23865
	,g23816,g23764,I22692,I22539,I22046,I22422,I22499,I22461
	,I21959,g22646,I22512,I22458,g22136,I22000,I22380,g22667
	,I22571,g23267,I22028,I22488,g22137,I21969,g22138,I22425
	,g22682,I22467,I22444,I22525,I21766,I21849,I22400,I22464
	,I22542,I22366,I22502,I22331,I22419,I21860,I21784,g25575
	,g22585,I21477,I21483,I23163,g24024,g24059,g24045,g24052
	,g24074,g24031,I22619,g24038,I21297,g24148,g24150,I21734
	,g25576,g22531,I21480,I26523,g24115,I22583,g24101,g24093
	,g24086,g24079,g24108,g24137,g24130,g24126,g24119,g24075
	,g24112,g24133,g24097,g24090,g24105,I22114,g24067,g24060
	,g24025,g24032,I22640,g24053,g24046,g24039,g24127,g24120
	,g24098,g24134,g24106,g24083,I22131,g24113,g24076,I23162
	,g24019,g24055,g24048,I22128,g24069,g24062,g24034,g24041
	,I21288,I21291,I22622,g24088,g24095,g24103,g24124,g24081
	,g24117,g24110,g24131,g25577,g23825,g24107,g24100,g24092
	,I22564,g24078,g24129,g24136,g24122,g24085,g24058,g24029
	,g24036,g24022,g24065,g24043,I22580,g24072,g24077,g24099
	,g24121,g24135,g24114,g24128,I22547,g24091,g24084,g24149
	,I21744,g24145,g24146,I21787,g24044,g24037,g24030,g24023
	,I22601,g24051,g24073,g24066,g24102,g24094,g24138,g24087
	,g24080,g24109,g24116,I22604,g24123,g24147,I21769,g24070
	,g24049,g24042,I22153,g24056,g24027,g24020,g24063,g24071
	,I22561,g24028,g24064,g24057,g24050,g24021,g24035,I21294
	,g24061,g24033,g24068,g24026,I22111,g24047,g24040,g24054
	,I21285,I21300,I21486,g24111,g24089,g24082,I22096,g24118
	,g24125,g24132,g24096,g24104,g16920,g18911,g23691,g23690
	,g25030,g21898,g24658,g25069,g24710,g24664,g25058,g21329
	,g23606,g24618,g24748,g25108,g17141,g23658,g25041,g24669
	,g24721,g25559,g22687,g22642,g22833,g22400,g25470,g25449
	,g25367,g20100,g20127,g20086,g21340,g21326,g19127,g20041
	,g23187,g25077,g23755,g22157,g21434,g24703,g23724,g22450
	,g25095,g24499,g24967,g23799,g21300,g23389,g20028,g22899
	,g24723,g22622,g17010,g24763,g25389,g25492,g16228,g23372
	,g24962,g25551,g22831,g24673,g16960,g21896,I20130,g25385
	,g16677,g25005,g25022,g24532,g21299,g23646,I21100,g24004
	,g25309,g25432,g25955,g24559,g22990,g23497,g24980,g25100
	,g25101,g25119,g24993,g19666,I22944,g15932,g25526,g25916
	,g24959,g24976,g24803,g24979,g25116,g24991,g25098,g25099
	,g23533,g25136,g25007,g25135,g25154,g25023,g22589,g25089
	,g23484,g22623,g25466,g24931,g24941,g24517,g24915,I19707
	,g23498,g22329,g23131,g21352,g17487,g23998,g22624,g19644
	,g24923,g23873,g23857,g23872,g25152,g22864,g21693,g21677
	,g23203,g21673,g23020,g23170,g21685,g23084,g21665,g21689
	,g23041,g21681,g21669,g23085,g23019,g23060,g21697,g23189
	,g21661,I22289,I22286,g21269,g23725,g26783,g24553,g25949
	,g23775,g23901,g23837,g23921,g23471,g23056,g17088,g24743
	,g25530,g24761,g19694,g22139,g24503,g22489,g22848,g22686
	,g23564,g23572,g24682,g22590,I19719,g24012,g19128,g23396
	,g23754,g22982,g23025,g24650,g20133,g23439,g25491,g21369
	,g23404,I21976,I19927,g17221,g23989,g23008,g22862,g21358
	,g23451,I22972,I20781,g25122,g24643,g24698,g25923,g23201
	,g21291,g18898,g23357,g25130,g25042,g21228,g23387,g24977
	,g23373,g24600,g16216,g22834,g24634,g23188,g22849,g22992
	,g25181,g25113,g22710,g24504,g26153,g23006,g20271,g25057
	,g23474,g21463,g25543,g25900,g24660,g20150,g25094,I20116
	,g25261,g25078,g21280,g23774,g24657,g23386,g23415,g23165
	,g24645,g22515,g21281,g23397,g23407,I21992,g23682,g25902
	,g22149,g22165,g22752,g22637,g22835,g22633,g21459,g21343
	,g22851,g17325,g23540,g26122,g16300,g22316,g16709,g24945
	,g24016,g24961,g24839,g22145,g22632,g22900,g24523,g23349
	,g24983,I20951,g24507,g22929,g22518,g22525,g23991,g23166
	,g24646,g23416,g25536,g24773,g24717,g23083,g21429,g25978
	,g21356,g24704,g24467,g21364,g20236,g25341,g25004,g24990
	,g21555,g25941,g25815,g26083,g25400,g21338,g25429,g24775
	,g25498,g25988,g23379,g24764,g25522,g25450,g25503,g25323
	,g22447,g25435,g24749,g25050,g24439,g24005,I20221,g20175
	,g19263,g20516,g20114,g20136,g20154,I16780,g20069,I16779
	,g25473,g25349,g20200,g24724,g21559,I20187,g25789,g21512
	,I20165,g24791,g25975,g19200,g20189,g20219,g19050,g20436
	,g18957,g18918,g25834,g25426,g25300,g26340,g25439,g24001
	,g23996,g23990,g24015,g26183,I20203,g25514,g26685,g23777
	,g20056,g25467,g24960,g25929,g24722,g25936,g25476,g21036
	,g25275,g24702,g23581,g23554,g25396,g24765,g25039,g25156
	,g25157,g25025,g25170,g23532,g23513,g23618,g23577,g23657
	,g25137,g25120,g25121,g24994,g25008,g22872,g24750,g25024
	,g25138,g25139,g25009,g25155,g25006,g25117,g25134,g25118
	,g24992,g24978,g24963,g25082,g25097,g25081,g24496,g24500
	,g24746,g24699,I25534,g25502,g25368,g25564,g24896,g19371
	,g21290,g19375,g19367,g19361,g21278,g19353,g21297,g23428
	,g24732,g24825,I23711,g26235,g26078,g26085,g25881,g25884
	,g25337,g25872,g25874,g25495,g26077,g26120,g26097,g26119
	,g26050,g24573,g25967,g22650,g22711,g22850,g26782,g24406
	,g23531,g26049,g26608,g25083,g24675,g25382,g22490,g25407
	,g25321,g25976,g26021,g24935,g24747,g25816,g26715,g25962
	,g24357,g23619,g23553,g24875,g24498,g26087,g26095,g24813
	,g25938,g26382,g23514,g25942,g26645,g26086,g24002,g22143
	,g24009,g21386,I24400,g26147,g26165,g24474,g24463,g26020
	,g26605,g24551,g25940,g25802,g26023,g25966,g26518,g25969
	,g20161,g25876,g25879,g25875,g25943,g26323,g26548,g25932
	,g26815,g26089,I24128,g26823,g26830,g25892,g20371,g21350
	,g25935,g21509,I25028,g25945,g23551,g23997,g25804,g25852
	,g25818,g26752,g23475,g25788,g24774,g21603,g25990,g26208
	,I23118,g24719,g26096,g25833,g25880,g26780,g26869,g26145
	,g26121,g24453,g25063,g24630,g26666,g25801,g26054,g25521
	,g24786,g24762,g25501,g25247,g26162,g25565,g26146,g25987
	,g26575,g25446,g25447,g24391,g24676,g25317,g24700,g25832
	,g26093,g24651,g24745,g24674,g26686,g26625,g25871,g26255
	,g26209,g26714,g26667,g21997,g21770,g22881,g21798,g21948
	,g21782,g21905,g21763,g21967,g21721,g25374,g21952,g21780
	,g21758,g21839,g21757,g21747,g21971,g22085,g21951,g21883
	,g21819,g21991,g21756,g21850,g22135,g21910,g21704,g21838
	,g22017,g21911,g21936,g21882,g22049,g21737,g21862,g21722
	,g21822,g22086,g21928,g22904,I24674,g24897,g21788,g21992
	,g22125,g21725,g22028,g22054,I24695,I24700,I24705,g23444
	,I24710,I24689,g21965,g21771,g25488,g22090,g22113,g22016
	,g21848,g21754,g22980,I24684,g21805,g22108,g22040,g21736
	,g22000,g21814,g21781,g21970,g22189,g25578,g21720,g21873
	,g21922,g21761,g21918,g21945,g21772,g21760,g21890,g23481
	,I27504,I27509,I27514,I26531,I27533,g22026,g23480,I24675
	,I24680,I24685,I24690,I24699,g21759,g21907,g21876,g21940
	,g22102,g24577,g24705,g21818,g22117,g22119,g21776,g22122
	,g21785,g21762,g21718,g21859,g22207,g21740,g21878,g22114
	,g22096,g22053,g21874,g21953,g22159,g25581,g21854,g21913
	,g22087,g23430,I27518,g22129,g21925,g22097,g22093,g24264
	,g21717,g21929,g21946,g22037,g21885,g23457,I24694,g21926
	,g21823,g21748,g24363,g22115,g21920,g25411,g22101,g21703
	,g22032,g22107,g21813,g25459,g22044,g21933,g22120,g22118
	,g23445,I27523,g22001,g21860,g22077,g24965,g21984,g22062
	,g23495,I27538,g21855,g21942,g21800,g22056,g21732,g22109
	,g22100,g22116,g21974,g22123,g21705,g21944,g22038,g21861
	,g22075,g22095,g21831,g21982,g21724,g22065,g21939,g22033
	,g21856,g22069,g22091,g21976,g22098,g22082,g21988,g21881
	,g21993,g21916,g22051,g22103,g22039,g22009,g21858,g21867
	,g22034,g22048,g22092,g21707,g22058,g25507,g21733,g21738
	,g21957,g22063,g21744,g22036,g21789,g21774,g24858,g21750
	,g21709,g21784,g21723,g21719,g21959,g21841,g22134,g22927
	,g24018,g21842,g21739,g21943,g25479,g21791,g21934,g21710
	,g22928,g21821,g21802,g22019,g25518,g22104,g22124,g21773
	,g21729,g22020,g21915,g23511,g21708,g22047,g24212,g21716
	,g21803,g21792,g21830,g21713,g21964,g21909,g21875,g22905
	,g21866,g23458,g21999,g25408,g21769,g21960,g21954,g21947
	,g22066,g21755,g21764,g21958,g21935,g22008,g22079,g21811
	,g21828,g21810,g21985,g21816,g21746,g22131,g22121,g21962
	,g22105,g21938,g21931,g22052,g21730,g21846,g22126,g21845
	,g21779,g22112,g21700,g22073,g21783,g21977,g22006,g21968
	,g21969,g21972,g21715,g22060,g21870,g21863,g21827,g21840
	,g21966,g25453,g21787,g21888,g22024,g21832,g21752,g21731
	,g22023,g21955,g21833,g21824,g21793,g21871,g21912,g21903
	,g21950,g21829,g22074,g21790,g22089,g22080,g21853,g24908
	,g21834,g21986,g21837,g21843,g22041,g21844,g22005,g22132
	,g22018,g21921,g21836,g21919,g21741,g22010,g21786,g21889
	,g21923,g22011,g22002,g22127,g22151,g22007,g21864,g21869
	,g22111,g21701,g21927,g24887,g21820,g21726,g22031,g22081
	,g25482,g22012,g22015,g22021,g21987,g21937,g21908,g22022
	,g21826,g22133,g22059,g21765,g21906,g25328,g22014,g24653
	,g21699,g21963,g21872,g25010,g22128,g22055,g21849,g22070
	,g22042,g21825,g21981,g25417,g21998,g21809,g21702,g22071
	,g21851,g21806,g22004,g21978,g21835,g22088,g22130,g21975
	,g21914,g23494,g21961,g21877,g21753,g22027,g22110,g22003
	,g24881,g21742,g21706,g21857,g21865,g21917,g21880,g21797
	,g21973,g22029,g22013,g21904,g22094,g21807,g21766,g21995
	,g21775,g21728,g24843,g21884,g21799,g24213,g22035,g21956
	,g21949,g22043,g21794,g22078,g21902,g21734,g21980,g22106
	,g21743,g22076,g21847,g21868,g21983,g21887,g21777,g22064
	,g21767,g21714,g22061,g21795,g22057,g21886,g21879,g21808
	,g21711,g21812,g22067,g21817,g21932,g22050,g22025,g22072
	,g21852,g21979,g21712,g22084,g21815,g21990,g21930,g22083
	,g21735,g21996,g21751,g21989,g22045,g21994,g22046,g21778
	,g21749,g21796,g22068,g21801,g22030,g21941,g21804,g21768
	,g21745,g22099,g21924,g22202,g22409,g23320,g23232,g23395
	,g23263,g23427,g23361,g23299,g22360,g22182,g23414,g23347
	,g23362,g23322,g22658,g24362,g23385,g22721,g23450,g23277
	,g22683,g23359,g23403,g22647,g23360,g23394,g23321,g22763
	,g23426,g23555,g22194,g22300,g22173,g22220,g22210,g23534
	,g23384,g23582,g23378,g23228,g23356,g23249,g23274,g23517
	,g23340,g23242,g23502,g23243,g23339,g23250,g23376,g23377
	,g23355,g23388,g23291,g23273,g23539,g23312,g23585,g23518
	,g23313,g23559,g23260,g23259,g23057,g23429,g22868,g22989
	,g22856,g22999,g23000,g23338,g22884,g23354,g23058,g23059
	,g22979,g23029,g23138,g23030,g23016,g22906,g23017,g22907
	,g23448,g23945,g23509,g23607,g23422,g23493,g24013,g23568
	,g23569,g23965,g23526,g23527,g23546,g23547,g23698,g23434
	,g23608,g23609,g23460,g23459,g23880,g23896,g23897,g22199
	,g23847,g23821,g23863,g23983,g23992,g23936,g22179,g22223
	,g22180,g23946,g23947,g23848,g23935,g23914,g23864,g23984
	,g22214,g23985,g23966,g23967,g23879,g22170,I21934,g23233
	,g23264,g23253,g23279,g23301,I22031,g23323,g23128,g22830
	,g23046,g23152,g23021,g22847,g23278,g23300,g22936,g23061
	,g23004,g23005,g22898,g22981,g23022,g22935,g23086,g23026
	,g23027,g22988,g22998,g23014,g23417,g23015,g23335,g22841
	,g23111,g22975,g22867,g22855,g22987,g23028,g22997,g22926
	,g23305,g22882,g22883,g23248,g23516,g23351,g23237,g23216
	,g23306,g23487,g23307,g23257,g23226,g23290,g23227,g23272
	,g23247,g23500,g23538,g23501,g23238,g23352,g23558,g23289
	,g23336,g23353,g23337,g23375,g23258,g22455,g22495,g22330
	,g22528,g22317,g22192,g22635,g22593,g22542,g23001,g22493
	,g23018,g22543,g22341,g22456,g22526,g22338,g22339,g22520
	,g22227,g22358,g22519,g22305,g23031,g22494,g22144,g23768
	,g23787,g23904,g23922,g22153,g23838,g23839,g23923,g23888
	,g23858,g23767,g23903,g23788,g23812,g22146,g22147,g23813
	,g23874,g23749,g23875,g23938,g22176,g22166,g23887,g23924
	,g23504,g23999,g23452,g23390,g23408,g23443,g23503,g23520
	,g23902,g23521,g23398,g23519,g23476,g23477,g23589,g23418
	,g23419,g23488,g23489,g23886,I21922,I21810,g23944,g22198
	,g23929,g23820,g23912,g23862,g23982,g23913,g22213,g23964
	,g23930,g23877,g23819,g23943,g22178,g22168,g22169,g23895
	,g22156,g23861,g23794,g23962,g23963,g23842,g23878,g23843
	,g23433,g23928,g23508,g23492,g23565,g23479,g23410,g23942
	,g24010,g23446,g23447,g23421,g23507,g23566,g23567,g23665
	,g23524,g23544,g23525,g23545,g22865,g22985,g23011,g23302
	,g23282,g22995,g22840,g23066,g22974,g22922,g22854,g22866
	,g22986,g23012,g23406,g22996,g23013,g22903,g22758,g22973
	,g23245,g23350,g23303,g23283,g23537,g23236,g23222,g23334
	,g23486,g23256,g23196,g23246,g23473,g23221,g23332,g23515
	,g23235,g23214,g23333,g23304,g23284,g23215,g23485,g23270
	,g23271,g23499,g23925,g23505,g23522,g23409,g23905,g23542
	,g23523,g23543,g23478,g23431,g23456,g23490,g23420,g23629
	,g23491,g23506,g23541,g24003,g23399,g23432,g23793,g23961
	,g23769,g23840,g22148,g23841,g23814,g23815,g23876,g23894
	,g23860,g23859,g23926,g22197,g23927,g23940,g23906,g23941
	,g23907,g23939,g23893,g22154,g23792,g22177,g22167,g22155
	,g22201,g23995,g22224,g23881,g23952,g23953,g22303,g23937
	,g23993,g23916,g23969,g23987,g23898,g23899,g22181,g23849
	,g23882,g23915,g22200,g24000,g22215,g23994,g23970,g23868
	,g23869,g23988,g23548,g23549,g23449,g23647,g23482,g23483
	,g23510,g23986,g23968,g24017,g23648,g23649,g23435,g23732
	,g23570,g23610,g23571,g23528,g23461,g23611,g24408,g26844
	,g25979,g24374,I21978,I22946,I21994,I22974,g24276,g24277
	,g25613,g25603,g25604,g25607,g25606,g25736,I22710,g24345
	,g24214,g24216,g25669,g25668,g26127,g24273,g24334,g24209
	,g24349,g24253,g24252,g24352,g25636,g21175,g24348,I22267
	,g24344,g25684,g26895,g24246,g24244,g25621,g24210,g24235
	,g25926,g25928,g25619,g24340,g25656,I21002,I20999,g24265
	,I20985,I20982,g25627,g25750,g26917,g24433,g24337,g24338
	,I21019,g24258,g24251,g24250,g26924,g24259,g24255,I22892
	,g24239,g24335,I22965,g26922,g24271,g24353,g24354,I21993
	,g24282,g24281,g24237,g24249,g25734,g25655,g24270,g26288
	,g24206,g24205,g24351,g26914,g22150,g26273,g25682,g25748
	,g25749,g25625,g19699,I24704,g24272,g25600,g25601,g26915
	,g24444,I22899,g26158,I22211,g24275,g25721,g24204,g25635
	,g24248,g25763,g24243,g24245,g25654,g24242,I20867,I20870
	,g25628,g24260,g25638,g24262,g25720,g25747,g24460,g24926
	,g25580,g24278,g26923,g25608,g25612,g24266,g25639,g20695
	,g24261,I21033,I21036,g19458,g24267,I22822,I21977,g24208
	,g24207,g25617,g25618,g25605,g24269,g24268,g24200,g24203
	,g24347,g26101,g26233,g25670,g24236,g24336,g18940,g24233
	,g24234,g25667,g24471,g24211,g24341,g24342,g24232,g24201
	,g25602,g25634,I22753,g25922,g25924,g25611,g25764,I22683
	,g25722,I20819,I20816,g24215,g24799,g25733,I27528,I24709
	,g24346,g25681,I22009,g23191,I23324,I23303,I23312,I23318
	,I23300,I23315,I23306,I23309,I23321,g25761,g24578,g24782
	,g24447,I24679,g25610,g25708,I20233,g24263,g24575,g26272
	,g18926,g25609,g25630,g24247,g25719,g24231,I22799,g26310
	,g25965,g24497,g25615,g26916,I19671,I19674,I22945,g26205
	,g26230,g26921,g26615,g26702,g26682,g26765,g21366,I22792
	,g24350,I20753,I20750,g26679,g19720,I20861,I20864,g24457
	,I22717,g25629,I20957,I20954,g26655,g26803,g26758,g26732
	,I20650,I20647,g24202,g25705,I22124,g24355,g25626,g24468
	,g25835,g25762,g25579,g24343,g25867,g25735,g25706,g24274
	,I21831,I22470,I22589,I22240,I22275,I22264,g26731,g24574
	,g24591,g25906,g25683,g25707,I20747,I20744,g25637,g25653
	,g24339,I20321,I20318,g23708,g23599,g23675,g23828,g23121
	,g22689,g22876,g22942,g22670,g23314,g23076,g23639,g23293
	,g23148,g23958,g23742,g23802,g22885,g22908,g26229,g22941
	,g26311,I21930,I22302,I21911,I22316,I22327,I22353,I21918
	,I22343,g25970,g26251,g26324,g23266,g25959,I22844,g22516
	,g22668,g26160,g26104,g24478,g26177,g22661,g25991,g22853
	,g22688,g26091,g26254,g26291,g25957,g22715,g26285,g26253
	,g25981,I22929,I22760,g25836,g25877,g26204,g26176,g26286
	,g26820,g26250,g22852,g22713,g26124,g26249,g25819,g22921
	,g26303,g26157,g22757,g25972,g26207,g26156,g26100,g26090
	,g26154,g26341,g24554,g25964,I22864,g22984,g26252,g26845
	,g26684,g26713,g26711,g26635,g25951,g23195,g26103,I20188
	,I20222,g26179,g26611,g22487,g26102,g25946,g26178,g25925
	,g25927,g24797,g24514,g24508,g24494,g26681,I22871,g26231
	,g22651,g25904,g26387,g27160,g24997,g25026,g24984,g24890
	,g24936,g24619,g27268,g26289,g24841,g26799,g26720,g26654
	,g26672,I22149,g26743,I22936,g27255,g22712,g26778,g23210
	,g22666,g27249,g22839,g26631,g27263,I20166,I20204,g27456
	,g23254,I24558,g26683,g22940,g27242,g24853,g24821,g24840
	,g24907,g27269,g26302,g26777,g26812,g26792,g26754,g26693
	,g26680,g26614,g23956,I21941,g22405,g22994,g22756,g22714
	,I22143,g26808,g26271,g27378,g26275,g26290,I22973,g23010
	,I20189,I22880,g26710,g26788,g26736,g26632,g14677,g23265
	,I22280,I22830,g22643,g22755,g22754,I21838,I22852,g25885
	,I20223,g25766,g26709,g24546,g25878,g25868,g27254,g27275
	,g26776,g26700,g26769,g26804,g26744,g27264,g26784,g26701
	,g26724,g24817,g24420,I22912,g23218,g26277,g22837,g26300
	,g26234,g22874,g26338,g25980,g26309,g27533,g25992,g26203
	,g25971,g26352,g25909,g25993,g22875,g27820,g25545,g27484
	,g23281,g22836,g25930,g22638,g25888,g26572,g25973,g26514
	,g22838,g26267,I22298,g27233,g26298,g27566,g22902,g26128
	,g26159,g26247,g26276,g26544,g27575,g27965,I25750,g27243
	,g26270,g24964,g26051,g27543,g27038,I20167,g26296,g27663
	,g26024,g26181,g26232,g26098,g26123,I20205,g26180,g27556
	,g27679,g25982,g27239,g27509,g27147,g26346,g26125,g26299
	,g27584,g26161,g26297,g26155,g26126,g25222,g25983,g25963
	,g26268,g26330,g26129,g26206,g24879,g24919,g24854,g27565
	,g27415,g25883,g26284,g27592,g27179,g27506,g27453,g26092
	,g26609,g26598,g26628,g26607,g25539,g25937,g27705,g24583
	,g24609,g27426,g24502,g27524,g27232,g26656,g26649,g26653
	,g27306,g24506,g27133,g26512,g27226,g27554,g27583,g27629
	,g27145,g27544,g27487,g26361,g26386,g26392,g27403,g26359
	,g27555,g26377,g27429,g26634,g26602,g25895,g25910,g27567
	,I22958,g27237,g27238,g27182,g27020,g27150,g26396,g26422
	,I23119,g27821,g27670,g26349,g25773,g27574,g27015,g26972
	,g27205,g27295,g27693,g27991,I23120,g27573,g27687,g27245
	,g27317,g26745,g26182,g24638,g22228,g22550,g24627,g22722
	,g22594,I23348,I23378,g25282,g25183,g25283,g25274,g25542
	,g25208,g25209,g24996,g25193,g25340,g24981,g24770,g25556
	,g25169,g25557,g25243,g25307,g25550,g25196,I24434,g25211
	,g25226,g25562,g25227,g25534,g25388,g25262,g24966,g25535
	,g25541,g25263,g25399,g24995,g25184,g25348,g25438,g25194
	,g24756,g25195,g24982,g25308,g25224,g25529,g25316,g25299
	,g25245,g25549,g25011,g25212,g25182,g25356,I23366,I23387
	,I23360,g26866,I23327,I23375,I23357,I23333,I23354,I23399
	,I23336,I23363,I23330,I23381,I23384,I23369,I23393,g24718
	,I23998,I24008,I24022,I24041,g25540,g24383,I24191,I24215
	,I24078,I23342,I23372,I23396,I23351,I23390,I23339,I23345
	,I24089,I24228,I24038,I24060,g24744,g25573,I23756,g26879
	,g24641,I26742,g25574,g26363,g25568,I23755,g25571,I24781
	,g26878,g24715,g25572,g25570,g25569,g25567,g20050,I25736
	,g22536,g24946,g24904,g25331,g26721,g26785,g26766,g26755
	,g26789,g26733,g26690,g24794,g24777,g25187,g24729,g25201
	,g25091,g20653,g24884,g25045,g25462,g27327,g27332,g24788
	,g24865,g27086,g27119,g23154,g23172,g23088,g23462,g23363
	,g22319,g22399,g22537,g25104,g24864,g27097,g25179,I22755
	,I22794,I22719,I22824,I22801,I22685,I22712,g24892,g24706
	,g22517,g22523,g27083,I23985,g25059,g27085,g22923,g24968
	,g25173,g25238,g27571,I23600,g20558,g25125,g24725,g25112
	,g26703,g26770,g26737,g25371,g24642,g21177,g27281,g25420
	,g20900,g25531,g20655,g25110,I22793,I22177,I22180,g25164
	,g25061,g25165,g24716,g23786,g18882,g25093,g24476,g24712
	,I22800,g24998,g25537,g25217,I22886,I22889,g26344,g25994
	,g25485,g19862,g24602,g24622,g24672,g24663,g24708,g24846
	,g27323,g24707,g24624,g22513,g22488,g24679,g26256,g25908
	,g24159,g24155,g24154,g24157,g24152,g24158,g24156,g24153
	,g24160,g24818,g22698,g25510,g25012,g24727,g24637,g25126
	,g26212,g25907,g24666,g20764,I22684,g25127,g25033,g25106
	,g27283,g25779,g25014,g25166,g25071,g25040,g26894,g24668
	,g24635,I22785,I22788,g25056,g25147,g25068,g24769,g25414
	,g24654,g24849,g26899,g24755,g25076,g22663,g26673,I22823
	,g25088,g24647,g24681,I22745,I22748,g21293,g24900,g25163
	,g25087,g23810,g24709,I22557,I24787,g26694,g25148,g24726
	,g24536,g26186,g27050,g22514,g22448,g25043,g24861,g25456
	,I22894,I22967,I22901,g25150,g22539,g22535,g25290,g25107
	,g20902,g25105,g24772,g25149,g27140,g25377,g23032,I22900
	,g25031,g27120,g27098,g24644,g24914,g24835,g25192,g24855
	,g25086,g24822,g22681,g24656,g25132,I22966,g24754,I22893
	,g25151,g24680,g24728,g25054,g21282,g25178,g21246,g25624
	,I24784,g21271,I23585,g27290,g25129,g25128,I22989,I23969
	,g24684,g25079,I25356,g24812,g28570,g26130,g24558,g24552
	,g27230,g25931,I22711,g25622,g27300,g27292,g27563,g27340
	,g25633,g22357,g22522,g23162,g27293,g28089,g25894,g26912
	,g25921,g26094,g25915,g26084,g26898,g28088,g22521,g25067
	,g23721,g25084,g27596,g28086,g26334,g26342,g24880,g28090
	,g25103,g27333,g24584,g24547,g28084,g27329,g27590,g25124
	,g25950,g25954,g23751,g27633,g22545,g22540,g26822,g19854
	,g22332,g24566,g23184,g24254,I22938,I22846,I22873,I22866
	,I22931,g19782,g24678,g26759,g27324,g26927,g26933,g27301
	,g28045,g26725,g19764,g26934,g22957,g22626,g26328,g26327
	,g27305,g22491,g22524,g19792,g24652,g28085,I22754,g25423
	,g24238,g27326,g25123,g25143,g26712,g26749,g26750,g26779
	,g28083,g24544,g24661,g26931,g26932,g25085,g28087,g22976
	,g27561,g26930,g27314,g27304,g26081,g25882,g25899,g25159
	,g28369,g27350,g25614,g27289,g25947,g25944,g27562,g26897
	,g26919,g26929,g26928,I22865,g25631,g26896,I22718,g26793
	,g27551,g27589,g27579,g25102,g27569,I22762,g25142,I26296
	,I22930,g23244,g22546,g23252,g23230,g23219,g22541,g23202
	,g22592,g24385,g24389,g24404,g24397,g24373,g24384,g24388
	,g24361,g24396,g24372,g25210,g25244,g25225,g25080,g25197
	,g24648,g25213,g25032,g24623,g25230,g24527,g24534,g24525
	,g24516,g24526,g24540,g24535,g24560,g24571,g24548,g24568
	,g24524,g24533,g24515,g24505,g24509,g24522,g24636,g25264
	,g25246,g25228,g25044,g25013,g25060,g28238,g27351,g27377
	,g26080,g26805,g28113,g28307,g27363,g27723,g28304,I22845
	,g27208,g27654,g28315,g28612,g27276,g28352,g27394,g27331
	,g28311,g28192,I22761,g28630,g28554,g28587,g25948,g25952
	,g27313,g27325,g27667,g25939,g28235,g28669,g27256,g25848
	,g27303,g27684,g27692,g28541,g28642,g27302,g27311,g27492
	,g27676,g27316,g27328,g28555,g28569,g27315,g28601,I22921
	,g27280,g27578,g27581,g28257,g27336,g27342,g27235,g28666
	,g27591,I22872,g27257,g27240,g27677,g27046,g25887,g27572
	,g27279,I22937,I25530,g28330,g27570,g27284,g27330,g27334
	,g27312,g28258,g28706,g27560,g28247,g28602,g28333,g28248
	,g27699,g28620,g27285,g28645,g26826,g25870,g25901,g26821
	,g27710,g27341,g28919,g23687,g28627,g27616,g26633,g28346
	,g27018,I26638,g28689,g27974,g27580,g27335,g28686,g24620
	,g28663,g28318,g27970,g27014,g28269,g28586,g25865,g27349
	,g28617,g23771,g24279,g28299,g27528,g27099,g27158,g27184
	,g28227,g28648,g28500,g28193,g27087,g28108,g28294,g28813
	,g23975,g23198,g25873,g25905,g26828,g23796,I26925,g27286
	,g27294,g27277,g27515,g27059,g27685,g28210,g28608,g28118
	,g25956,g25958,g28215,g28144,g28154,g26335,g26329,g29172
	,g27463,g27041,g27017,g27552,g27291,g26343,g26348,g28441
	,g26099,g28159,g28324,g28339,g27646,g27717,g27247,g28151
	,g28812,g27597,g28117,g28321,g28219,g28633,g24314,g24300
	,g25141,g24291,g24326,g24327,g24191,g24299,g24333,g24288
	,g24189,g25504,g24289,g24306,I25612,I25613,g24226,I25359
	,g24190,g24287,I25219,g25640,g24194,g24324,g24301,g24197
	,g24218,g24286,g24298,g24329,g24293,g24186,g24308,g24230
	,g24323,g24316,g24319,g24229,g24561,g24220,g24187,g24193
	,g24188,g24312,g24227,g24302,g24295,g24292,g24228,g24322
	,g24195,g24330,g24222,g24309,g24304,g24283,g24224,g24196
	,g24297,g24221,g24320,g24290,g24285,g24332,g25694,g24303
	,I25327,g24313,g24307,g24219,g24294,g24223,g24311,g25693
	,g24225,g24217,g24199,g24310,g24296,g24198,g24317,g24325
	,g24305,g24284,g24331,g24321,g24315,g24328,g24192,I25242
	,g24318,g24893,g24866,g25064,g24920,g24911,g25051,g25027
	,g24869,g24850,g24836,g24819,g27008,g27511,g25250,g24490
	,g24366,g24377,g24407,g25563,g24365,g25538,g24386,g24356
	,g25544,g25558,g25528,g25552,g24426,g24376,g24438,g24418
	,g24419,g24424,g24364,g24425,g24375,g24428,g24429,g24405
	,g24452,g24431,g25553,g24367,g25523,g24358,g24359,g25546
	,g25547,g24379,g25554,g25566,g25555,g25560,g25525,g25561
	,g25533,g25548,g25452,g25326,g25409,g24394,g24360,g25517
	,g25410,g25286,g25287,g25480,g25231,g25481,g25370,g25451
	,g25140,g25324,g25506,g25325,g25214,g24368,g25185,g25524
	,g25266,g25267,g25288,g25289,g25158,g25171,g25198,g25232
	,g25369,g25505,g25248,g25249,g28677,g28451,g28456,g25688
	,g26424,I23986,I23601,I23586,I23970,g25752,g25677,g23575
	,g24933,g24972,I23971,g24943,g23823,g25019,g25731,g25744
	,g24958,g25021,g28077,I23587,g26940,g25742,g24989,g23824
	,g25641,g28043,g23800,g25741,I22576,g25701,g25002,g27858
	,g27800,g25679,g24942,g24934,g25650,g25651,g25759,g25758
	,g23761,g24917,g25661,g23809,g25757,g25662,g26939,g24688
	,g26515,g26616,g25730,g28078,g25698,g25697,g25592,g25649
	,g26545,g28578,g25755,g25595,g25599,g25648,g28076,g28075
	,g25710,g25695,g23762,g25678,g28518,g24924,g25770,g25821
	,g25532,g25739,g25740,g25594,g25712,g25711,g23746,g26865
	,g25791,g27907,g25745,g25777,g25729,g26574,g26657,g25223
	,g24518,g25724,g25728,g25690,g28070,g26938,g25691,g25660
	,g25726,g25727,g27265,g27614,g27251,g27594,g27975,g27088
	,g25642,g23440,g25700,g25357,g25702,g25703,g26603,g24918
	,g23870,g23613,g25665,g25664,g25672,g25716,g23685,g25003
	,g27600,g27259,g27246,g27588,g27971,g27084,g25207,g24510
	,g25666,g25676,g25674,g25675,g25689,g25769,g25805,g25715
	,g25713,g24957,g25717,g25723,g25714,g23653,g25658,g25381
	,g25737,g25048,g25709,g23616,g25671,g25725,g23552,g23715
	,g24916,g25663,I25845,g25685,g28073,g25673,g24951,g25696
	,g25049,g25800,g25856,g26337,g25038,I25907,g24906,g25645
	,g25646,g25425,g25597,g25657,g25659,g26546,g26636,g24974
	,g25746,g25644,g25643,I22816,I22819,g25784,g25839,g25743
	,g25593,g24944,g27585,g25020,g23760,g24975,g24932,g25756
	,I25586,g23656,g25686,g24925,g25751,g22171,g25018,g25591
	,g25062,g25753,g25760,g23003,g23655,g23651,I25594,g23745
	,g23576,g25778,g23776,g25754,g26872,g27601,g27260,g27092
	,g27984,g27266,g27615,g27990,g27101,g27595,g27252,g27089
	,g27976,g25647,g25699,g23529,I23602,g25527,g25704,I24445
	,I24448,g28071,g28072,g25738,g25596,g28074,g24950,g28591
	,I24117,g25598,g25785,g26573,g23650,g25687,g25732,g25718
	,g25652,g26484,g26398,g25680,g26873,g23231,g24485,g24537
	,g24541,g24491,g24872,g28544,g24905,g27634,g27270,I24497
	,I23671,I24455,I23680,I23684,I23694,I24474,I23688,g26485
	,g26516,I23949,g23719,g24988,g23780,g24973,g23617,g28534
	,g27662,g27598,g27648,I23987,g27994,g27112,I24383,g25632
	,g23747,g28564,g28545,g28536,g28056,g27958,g27962,g24567
	,g23748,g28613,g28577,g24621,g27576,g28549,g26944,I24334
	,I24331,g23781,g27102,g27093,g24601,g27019,g24929,g27025
	,g27028,g27742,I25190,g27779,g24631,g27091,g27983,I24414
	,g29293,g27100,g27989,g28165,g28581,g25960,g25623,g28592
	,g26918,g24549,g28712,g28697,g28695,g28679,g28658,g22873
	,g22938,g28110,g28676,g28692,g28638,g28655,g22920,g22861
	,g28107,g28657,g28674,g28714,g28725,g29837,g28426,g27362
	,g28455,g28532,g28341,g28710,g28694,g28582,g26864,g28182
	,g28603,g28551,g29302,g29264,I23961,g27959,g27963,g26079
	,g26920,g26829,g26048,g26019,g24662,g27278,g27542,g27532
	,g27274,g24921,g28052,g25866,g29282,g29283,g28167,g28558
	,g24570,g24555,g29299,g25986,g25831,g26925,g29296,g27029
	,g27034,g26833,g28448,g29273,g28055,g29078,g27886,g27837
	,g26855,g29265,g29266,g28044,g29295,g27937,I22922,g24677
	,g29301,g29300,g28595,g29306,g29307,g28137,g29272,g26301
	,g28574,g26926,g28060,g29284,g26913,g26088,g28580,g29224
	,g26274,g28576,g24576,g29270,g28548,g28605,g28054,g28204
	,g28353,g28513,g26838,g29294,g28526,g28051,g25850,g27957
	,g27932,g29271,g29305,g29261,g26839,g29308,g28152,g28561
	,g28594,g28525,g29267,g26818,g29190,g29288,g26847,g28546
	,g28058,g28607,g28596,g26287,g26279,g28517,g26846,g28565
	,g29290,g29287,g28566,g26854,g26294,g28047,g26292,g28560
	,g29289,g29281,g26849,g28050,g28049,g26848,g28046,g28562
	,g28589,g26304,g25782,g25775,g26853,g29260,g26312,g25768
	,g28479,g26257,g29259,g26842,g28625,g29258,g28614,g26858
	,g27224,I24363,g28198,g27250,g27016,g27393,g29643,g27964
	,g27968,g27612,g28533,g29933,g29475,I22923,g24949,g27024
	,g28573,g28174,g28653,g28538,g24912,g28160,g28325,I24461
	,g30184,g24939,I23978,g29196,g28597,I26989,g28527,g27026
	,g28431,g28164,g28504,I23917,g29325,g28279,I24438,g29745
	,g28368,g28370,g27036,g27043,g27035,g27030,g24564,g28444
	,g29477,g27231,g27258,g29319,g30173,g28314,g28285,g28672
	,g28598,g29114,g28237,g25838,I25562,g25783,g25869,g28180
	,I26710,I27492,g28119,I25221,g26827,g26831,g26832,g26837
	,g25790,g25820,I25146,I25161,g25837,g26836,g26841,I25244
	,g26082,g26364,I24759,I24839,I25677,I25220,g26483,g26874
	,g26365,g24891,g27366,g26604,g26547,g27027,g26976,g27400
	,g26541,g27703,g27771,g27368,g26381,g25240,g27875,g27954
	,g27770,g27823,g25765,g28796,g28966,g27704,g27354,g25774
	,g26511,g27926,g24808,g28843,g28874,g28837,g28903,g27722
	,g25260,g27927,g29248,g25780,g24380,g26166,g26148,g25180
	,g27382,g25380,g26819,g27982,g28765,g28935,g25296,g26860
	,g25241,g26190,g26213,g26308,g27826,g26630,g26652,g28871
	,g28942,g26358,g26394,g26399,g27924,g24759,g26380,g26379
	,g26357,g26395,g26391,g26389,g27647,g26857,g27828,g24417
	,g27829,g26612,g28946,g28994,g29131,g29134,g26856,g26852
	,g29225,g25298,g26871,g27010,g27879,I26667,g25772,g27337
	,g23684,g28236,g28245,g27721,g26863,g25767,g28867,g28793
	,g29057,g29060,I25908,I25909,g26513,g26650,g26542,g26651
	,g26670,g26671,g27599,I26960,I27409,I27381,I27429,I27364
	,I26972,I27349,I26948,g27356,g27338,g26689,g26360,g27732
	,g26517,g27735,I25846,I25847,g26571,g26543,g27733,g26486
	,g26390,g25272,g26393,g26347,g27768,g27364,g26258,g26356
	,g26325,g27343,g26613,g25917,g25221,g26362,g26378,g27966
	,g26200,g26241,g26313,g26423,I25692,g27353,g27659,g25781
	,g26861,g27731,g26388,g25206,g25513,g27516,I24278,I24281
	,I25683,I25695,g27960,g27007,g26261,g26223,g25786,g27969
	,g27720,g26339,g26397,g26487,g29170,g29152,g29130,g28713
	,g26351,g25297,g26244,g26281,g26226,g26264,g26753,g26719
	,g26336,g28907,g28840,g29097,g29094,g29092,g29056,g29128
	,g28678,g28696,g29093,g29129,g29151,g23453,g25424,I25680
	,g25465,g24369,g29227,g26259,g27369,I24237,I25243,g24802
	,I25786,I25779,I25790,g27730,I25689,g26306,g26350,g26295
	,g26307,g26345,g26280,g26610,g26629,g27697,g27696,g30125
	,g27673,g27674,g27288,g27287,g30110,g30135,g30066,g30099
	,g27683,g27682,g28178,g27665,g27666,g30094,g30084,g27299
	,g27298,g30095,g27691,g27690,g27310,g27309,g30121,g30086
	,g30122,g30133,g30158,g27660,g27766,g27479,g29049,g29046
	,g28857,g28920,g27652,g27827,g27772,I23950,g27877,g27973
	,g27367,g29275,I24384,g27352,g26993,g27345,g27012,g26800
	,g27734,g28911,g28973,g28783,g28758,I24415,g27825,g25996
	,g27355,g28547,g28524,g28535,g28563,g27381,g28537,g28567
	,g28550,g28583,g25911,g26606,g26236,g26218,g26195,g26171
	,I24416,g28268,g28246,g28284,g28256,g28824,g28892,g27769
	,g27344,g29115,g29080,g29045,g28675,g26187,g28656,g29079
	,g29014,g29044,g28208,g27379,g27878,g28121,g28127,g27499
	,g25168,I26654,g28134,I24385,g28149,I27192,g24952,g27063
	,g24483,g25284,g24489,g24481,g24477,g25265,g24466,g25322
	,g26326,g25849,g25893,g25886,g25830,g28830,g28864,g29242
	,I23951,g25984,g29247,g29246,g25995,g29230,g26781,g29243
	,g29223,g28853,g28780,g29255,g29241,g28736,g28755,g28048
	,g28931,g28987,g29118,g29121,g29253,g23778,g29226,g29235
	,g30049,g29359,g28255,g28265,g29240,I26004,g29245,g28927
	,g28861,g28877,g28914,g29229,g26278,g29250,g28132,g28900
	,g28962,g29660,g28885,g28820,g29015,g29018,g28786,g28955
	,g24240,g29507,g29254,g30334,g25985,g26025,g25953,g26052
	,g26293,g24241,g29025,g28977,g29154,g29157,g30671,g29378
	,g24257,g29251,g29001,g28950,g29177,g29171,g28726,g29153
	,I23962,g29149,g29081,g29116,g28693,g28711,g29117,g29169
	,g29150,g29513,g29228,g28211,g29333,g29252,g29244,g29834
	,g24256,g28135,I23963,g29249,g29583,g30089,g30126,g30137
	,g30161,g28442,g28626,g30078,g30112,g30124,g30149,g30111
	,g30098,g28185,g28440,g28616,g30109,g30075,g30145,g30120
	,g30108,g30051,g30083,g30118,g28301,g28415,g28183,g28171
	,g29324,g30107,g30064,g30131,g30096,g30139,g30101,g30172
	,g30151,g30138,g31252,g29746,g25974,I24439,g29367,g29082
	,g29085,g28896,g28827,g26751,g29924,g29916,g29376,I24440
	,g26053,I23918,g28053,I23979,g29707,I24462,g30322,g29744
	,I28576,g29679,g29329,g28508,g29256,g26809,I24364,g29494
	,I24463,g26813,g29508,g30287,g31509,g30982,g29343,g31243
	,g28138,g29706,I24365,g30062,g29361,g30935,g29330,g29937
	,g26305,I23980,g30291,I28128,g29668,g31654,g29375,I23919
	,g28427,g28313,g31144,g29597,g28212,g28216,g29778,g29363
	,g30579,g29570,g29793,I26530,g27649,g27627,g28040,g28034
	,g28038,g28039,g28032,I26100,g28033,g28036,g28037,g26248
	,g26935,g25692,g25620,g27414,g27467,g27439,g27493,g26269
	,g26131,g26105,I27758,g29194,g28187,g29385,g26840,g27042
	,g27033,g26881,g26880,g26961,g26966,g26968,g26962,g26967
	,g26963,g28803,g26941,g27074,g27051,g27064,g29954,g28223
	,g27057,g26314,g26886,g27550,g29519,g25073,g27032,g28082
	,g26964,g29628,I25606,g26936,I25598,I24393,I24396,g26946
	,g27185,g29360,g28477,g27058,g29576,g28197,g30088,g30020
	,g30038,g30079,g29913,g29953,g28115,g26965,g28499,g26892
	,g29883,g27045,g29968,g26893,g28010,g28020,g27617,g27602
	,g27999,g26977,g26994,g27635,g29612,g28478,g26900,g26908
	,I25579,g26906,g28454,g26956,g27738,g27833,g27882,g27775
	,g26905,g29364,g26902,g27044,g28232,g28543,g27225,g28202
	,g27651,g28523,g26943,g26970,g29732,g30298,g26937,g25115
	,g29604,g28240,g26947,g29651,I24920,g26811,g26952,g26903
	,g26904,g30293,g28272,g28139,g26942,g26958,g26890,g26907
	,g26969,g28531,g26901,g26814,g27011,g28116,g27613,g26971
	,g26945,g26949,g26960,g29588,g29596,g26889,I25567,g26951
	,g26953,g26909,g26910,g27141,g28225,g26954,g26957,I26522
	,g28260,g28300,g28124,I26936,g26888,g26882,g26887,g26883
	,g27223,g29711,g30019,g30067,g29997,g30077,g29906,g29942
	,g27931,g25242,g28489,g28156,g28273,g26824,I26430,g30039
	,g30054,g30090,g30100,g30021,g29967,g27759,g27711,g27450
	,g26911,g26955,g29528,I25005,g28244,g27587,g27724,g27700
	,g26950,g26260,g26948,g29981,g29928,g26891,g27031,g29525
	,I25555,I26448,g27161,I25576,g29980,g30299,I25591,I25541
	,g28599,g26816,g29965,g29922,g29923,g30313,g29642,g26884
	,g29998,g30306,I25552,g26959,g26885,I25369,g27586,g29501
	,g29313,g29362,I25115,I25351,I25095,I25366,I25380,I25399
	,I25105,I25391,g25776,g25851,g30003,g24792,g27146,g28068
	,g30369,g28214,g28234,g28136,g28098,g29637,g30366,g29940
	,g28104,g27577,g29535,g28251,g28064,g28095,g27209,g29882
	,g29512,g27668,g27122,g30352,g28709,g27593,g28213,g30378
	,g29577,g28133,g29870,g29854,g29585,g29587,g28217,g30364
	,g29838,g28091,g29688,g29683,g28103,g28312,g29943,g28148
	,g29662,g27040,g30300,g29486,g29496,g30314,g30307,g29489
	,g25215,g28466,g28572,g29804,g29686,g29868,g29687,g29551
	,g29605,g28289,g29869,g28101,g30365,g27714,g27762,g29621
	,g28243,g29603,g27468,g27727,g27817,g27162,g29553,g29895
	,g28100,g28147,g29619,g28557,g28494,g30371,g29664,g28112
	,g30304,g30311,g28218,g29615,g28200,g29665,g26718,g27210
	,g28094,g29840,g28229,g27261,g28495,g28111,g28065,g28242
	,g29600,g29851,I26409,I26406,g29710,g28062,g29238,g28130
	,g27658,g27039,g30372,g28067,g28467,g29482,g29488,g29582
	,g29961,g29920,g28205,g27073,g28097,g30363,g25236,g29566
	,g29485,g29495,g29636,g27037,g27009,g28488,g27796,g27933
	,g27903,g27854,g29649,g29547,g30353,g30370,g30297,g29905
	,g29999,g29944,g30367,g28199,g29620,g29855,g28061,g28233
	,g30351,g29977,g29939,g30074,g29994,g30065,g30016,g28092
	,I26799,g27988,g29969,g30091,g29985,g30080,g27541,g27992
	,g29381,g29380,g29629,g29377,g29613,g27553,g31238,g25096
	,g29521,g29865,g29509,g29645,g28201,g28261,g29511,g24798
	,g29538,g27108,g27664,g29731,g30333,g29853,g28143,g29573
	,g27217,g29584,g27248,g27241,g29926,g29964,g28226,g31294
	,g29839,g29631,g27186,g29648,g28125,g29955,g30022,g30566
	,g30456,g31894,g29646,g29574,g27121,g29852,g29601,g30102
	,g30055,g30068,g30113,g29983,g30040,g29514,g27244,g29995
	,g30303,g29602,g29976,g30052,g29993,g30063,g29925,g29960
	,g29996,g29941,g27765,g29929,g29312,g29563,g29927,g29978
	,g27822,g27320,g29617,g27686,g30053,g30037,g30087,g30097
	,g30018,g29963,g29893,g30292,g28585,g29911,g29948,g27678
	,g29524,g29921,g30310,g29276,g29532,g29867,g29638,g29685
	,g30362,g25199,g31271,g30349,g29599,g30377,g30387,g29661
	,g29709,g30670,g30360,g30361,g29684,g29530,g30348,g29633
	,g29951,g29279,g31527,g29568,g29634,g30356,g29667,g30355
	,g29233,g30376,g30368,g29894,g30354,g29517,g29586,g32053
	,g32296,g30383,g29589,g30386,g29733,g30375,g29549,g29616
	,g29622,g30357,g30335,g32201,g31523,g29572,g31866,g27564
	,g29708,g29712,g30380,g30374,g30359,g30381,g29866,g27253
	,g31149,g31014,g29984,g30379,g31247,g27997,g29884,g29652
	,g25271,g29740,g29881,g29880,g30350,g31221,g30384,g24807
	,g29907,g27995,g30373,g29663,g32019,g31013,g29237,g29896
	,g30325,g31227,I28913,g27236,g30336,g29232,g27271,g24760
	,g29278,g29277,g25258,g31239,g31668,g29234,g27981,g29912
	,g29950,g30076,g30036,g30017,g30085,g29231,g30385,g30382
	,g30358,g30023,g29383,g29644,g29630,g30607,g30600,g32197
	,g29564,g31262,g30936,g30612,g30918,g29236,g29239,g31134
	,g30577,g31020,g30342,g31964,g29897,g32040,g31670,g32155
	,g30731,g30730,g31233,g31277,g31474,g31138,g31069,g31848
	,g31849,g31805,g31798,g31813,g31799,g31852,g31808,g31809
	,g31836,g31853,g31822,g31837,g31830,g31842,g31816,g31823
	,g31817,g31810,g31843,g31831,g31856,g31857,g31802,g31850
	,g31811,g31826,g31803,g31827,g31846,g31820,g31851,g31847
	,g31840,g31796,g31797,g31834,g31821,g31806,g31835,g31841
	,g31807,g31814,g31800,g31815,g31838,g31839,g31854,g31801
	,g31818,g31819,g31855,g31824,g31844,g31858,g31825,g31859
	,g31832,g31845,g31828,g31829,g31812,g31833,g31804,I27543
	,I28062,g29474,g27980,g27972,g26990,g27977,g26973,g27142
	,g27004,g26987,g27155,g27985,g27282,g28340,I27508,I27513
	,g28326,g28035,I27539,I27534,I27519,I27524,I27529,g27402
	,g28476,g28521,g27582,g26510,I27503,g28491,g28482,g29186
	,g31142,g31147,g29479,g28888,g28253,g28059,g30081,g31007
	,g29848,g31776,g29892,g29484,g28981,g28953,g26834,g29193
	,g28106,g31319,g31472,g29776,g31307,g28990,g28186,g28290
	,g28637,g30163,g28363,g28376,g28406,g28391,g28395,g28381
	,g28410,g28421,g29480,g29167,g29146,g29792,g30176,g27961
	,g31210,g29849,g29173,g29187,g29370,g26825,g28965,g28934
	,g29184,g29181,g28856,g28823,g26859,g30141,g26850,g28923
	,g28263,g27929,g31169,g26835,g31790,g31375,I26195,g28031
	,g28057,g29692,g28559,g28590,g29007,g28986,g25903,g29107
	,g29180,g29175,g29069,g29034,g28575,g28604,g27881,I26516
	,g30115,I27677,g31152,g29502,g31788,g26817,g29864,g28457
	,g28452,g31186,g28492,g28483,g28475,g28209,g28443,g29786
	,g29070,g29756,g29035,g29012,g28930,g29775,g30189,g26843
	,g29072,g29040,g28414,g27395,g27421,g27416,g27445,g31001
	,g29141,g29104,g27474,g27494,g27440,g27469,g28520,g28515
	,g29109,g29077,I26508,g29164,I26644,g29142,g31131,g31141
	,g30103,g28895,g28860,I26581,g28480,g28469,g29174,g29165
	,g29735,g31778,I29207,I26503,g25771,g30564,g28584,g28540
	,g28498,I26643,g28493,g26648,I29211,g27669,I26584,g30104
	,g29148,g31759,g29145,g29005,g29198,g29183,g29106,g29071
	,g28425,g26851,g27273,g31787,g31777,g25220,g26862,g26870
	,I25511,I25514,g28380,g28241,g28109,g28131,g28114,I27401
	,g28250,g28399,I26578,I28185,I28199,I27927,I28174,I27941
	,I27954,I27970,I28162,g28158,g28274,g28153,g31293,g29716
	,g29108,g29144,g28462,g28470,g28468,g29717,g29791,g30201
	,g28519,g28552,g29006,g29032,g28624,g29777,g29189,g29200
	,g25968,g28481,g30127,g25787,g29487,g28280,g28899,g28958
	,g29476,g28302,g29028,g30093,g28510,g28514,g29768,g30128
	,g31130,g31124,g29033,g28529,g28568,g29879,g28496,g28509
	,g29191,g29179,g28282,g28191,g28969,g28194,g28673,g29506
	,g31168,g29753,g30114,g30092,I29261,I29277,g29741,g29748
	,g29790,g29483,g29168,g29478,g29754,g27832,g29763,g31002
	,g31187,I29269,g28292,g27737,I29284,I29313,I29225,I29218
	,I28548,g29802,g28266,g28615,g28593,g30214,g29904,g28606
	,g28579,g29801,I29221,I29228,I29214,g29490,I28241,g28126
	,I25869,I25882,g26549,g26026,g26576,g26519,g26488,g25997
	,g26400,g26055,I29242,g28096,I29295,g31209,g31148,g31153
	,g28066,g28976,g31185,g31123,g31128,g30340,g30346,I29302
	,g30392,g31151,g28906,g28870,g30341,g31211,g28938,g30389
	,g31222,g28949,g28997,I27235,I27238,g29734,g28063,g29813
	,g25977,g30338,I29253,g29004,g29504,g30390,g28980,g31166
	,g28945,g28910,g29481,g28654,g28188,g29764,g32424,g30339
	,g28099,g31867,g25803,g25616,g28120,g30391,g31948,g32425
	,g32169,g32207,g32254,g31145,g31139,g31129,g32034,g33299
	,g33124,g25817,g28093,g28069,g31150,g31962,g33035,g30931
	,I29371,g32037,g31122,g31120,g28102,g28105,g31865,g25961
	,g32395,g31146,g31140,g33258,g31864,g30388,g32978,g30347
	,g31167,g30345,g32399,g30344,g33126,g31870,g26022,g33235
	,g25814,g25989,g32011,g32173,g31184,g33113,g32137,g31868
	,g32125,g32192,g31524,g32339,g31934,g31963,g33252,g32181
	,g32041,g32212,g32094,g32190,g32012,g32154,g32138,g32016
	,g32202,g28512,g28522,g28516,g29208,g29203,g29202,g28652
	,g28288,g28271,g28298,g28259,g28287,g28270,g28203,g28206
	,g28207,I26952,I26929,I28579,g29814,g29209,g32341,g31494
	,g31769,g31517,g29338,g31784,g31519,g32316,g31750,g31125
	,g31475,g32160,g31270,g32327,g31485,g31786,g31752,g29327
	,g31707,g31484,g31516,g31780,g29314,g29369,g29334,g31018
	,g31017,g29332,g31525,g32334,g31758,g32166,g31292,g31067
	,g31490,g30025,g29930,g29713,g29689,g29669,g29945,g29653
	,g29970,g29956,g29503,g29497,g28079,g29067,I28434,g30026
	,g30004,g29835,g29803,g29850,g29836,g28264,g29571,g29579
	,g29592,g29606,g26802,g30069,g30058,g31504,I26466,I26451
	,g26810,g28970,g28939,g29548,g32219,g29354,g29975,g29990
	,g29609,g29624,g29345,g30009,g30028,g28991,g28959,g30286
	,g29531,I26381,g29029,g28998,g30056,g30044,g29959,g29973
	,g30034,g30047,g29719,g29657,g28081,g32275,g32222,g31609
	,g27698,g28140,g29656,g29641,g32228,I26479,g27993,g28303
	,g31601,g28080,g29352,g27996,g30059,g30048,g28172,g28179
	,g32262,g29349,I26356,I26741,g28453,g29336,I28458,g29346
	,I26512,g32236,g29351,g29317,g29737,g29676,g29694,g29672
	,g28009,I27368,g29722,g29702,g29534,g29550,g29647,g29522
	,I25743,g29598,g29510,g29515,g29206,g29201,g29205,g29204
	,g29207,g27527,I26337,g32249,I27391,I26378,I26427,I26309
	,I27495,g29878,g29863,g29812,g29847,g29846,g29862,g29811
	,g29800,g32223,I26334,g29505,I26130,g30073,g29625,g29639
	,g27096,g27213,g28230,I29314,g31658,g27187,g27163,g27126
	,g29567,g29974,g29988,g30071,g30082,g30070,g30060,g28283
	,g30279,g29350,g30012,g28799,g28761,g28833,g28789,g28739
	,g28846,g28768,g28880,g29675,g29705,g30007,g30027,g30006
	,g29989,g29575,g31616,I29270,g31646,g31631,I29285,g27405
	,g29565,g32247,g28267,g29578,g28291,g29632,g29523,g29533
	,g29991,g30008,g30033,g30045,g30032,g30015,g30029,g30042
	,g32211,g29536,g29614,g29516,g29569,g28293,g30301,g32218
	,g31624,g31639,I29315,g29580,g29591,I29286,I27449,g29611
	,g29626,g29610,g29595,g32264,g30011,g30030,g30010,g29992
	,g28439,g28254,g28889,g28918,g28924,g28281,g29607,g29623
	,I29278,g29640,g29627,I29279,I29262,g30043,g30031,g29348
	,g29593,g29581,g30057,g30046,g30270,g29355,g29335,I28002
	,g30318,I28572,g29339,I28014,g31792,g31765,g31500,g31540
	,g29321,g31471,g31492,g31746,g31477,g29986,g31015,g31016
	,g31278,g31066,g31520,g31499,g31756,g31478,g29344,g31470
	,g31744,g32308,g31374,g30002,g31115,g31280,g31132,g31290
	,g31481,g32162,g31508,g31493,g31763,g31789,g31486,g31118
	,g31305,g31143,g31019,g27411,g27557,g27508,g27537,g27538
	,g27546,g27507,g27460,g27136,g27129,g27104,g27114,g27262
	,g27218,g27135,g27517,g27480,g27428,g27370,g27346,g27427
	,g27481,g27385,g32271,g27653,g27547,g27116,g27130,g27181
	,g27204,g29608,g29594,g30061,I26438,g27220,g27203,g27106
	,g27151,g27115,g27214,g27219,g27137,g27105,g27180,g27373
	,g27387,g27267,g27227,I30904,g27134,g27177,g27103,g27095
	,g27212,g27211,g27094,g27202,g27148,g27128,g27645,g27534
	,g30050,g29342,g27389,g27486,g27545,g27520,g27521,g27433
	,g27485,g27535,g27650,g27536,g27347,g27371,g27500,g27358
	,g27437,g27462,g32243,I29263,I29296,g29552,g27431,g27207
	,g27132,g27234,g27221,g27206,g27154,g27228,g27222,g27272
	,g27229,I29254,g27457,g27375,g27504,g27409,g27361,g27505
	,g27201,g27149,g27113,g27178,g27127,g27090,I26070,g27372
	,g27360,g27482,g27430,g27519,g27518,g27454,g27407,g27359
	,g27503,g29590,g27490,g27461,g27526,g27540,g27215,g27183
	,g27118,g27216,g27139,g27107,g27404,g27357,g27501,g27451
	,g27628,g27339,g27452,g27384,I26459,I29255,g32210,g27376
	,g27522,g27390,g27410,g27434,g27459,g32285,g32229,g27408
	,g27374,g27432,g27388,I29271,g27117,g27131,g27138,g27153
	,g28754,g32216,I26366,I26049,g27455,g27386,g27502,g27348
	,g27483,g27406,g27391,g27488,g27435,g27523,I26393,g32277
	,g29537,g29618,g29518,I29303,g27525,g27412,g27558,g27549
	,g27491,g27436,g27413,g27539,g27559,g27510,g32237,g32235
	,I29304,I26417,g27548,g27568,g27392,g27661,I26093,g32259
	,I29297,g27383,g32976,g32209,g32233,g32220,g32221,g29526
	,g29650,g29554,g32217,g29527,g29635,g29666,g29555,g32227
	,g32982,g32981,g33723,g33851,g32977,g27152,g32208,g31795
	,I29717,I29720,g30035,g33123,g32980,g33799,g32226,g33102
	,g33099,g33817,g33186,g33241,g33245,g33122,g33232,g33724
	,g27458,g33615,g32257,g27489,g33794,g32245,g27159,g32985
	,g31872,g33019,g33121,g33306,g33104,g32984,g33291,g33244
	,g33538,g33233,g33246,g32979,g33322,g33105,g33159,g30326
	,g28436,g28463,g29752,g29736,g29718,I28480,g27438,g30599
	,g30595,g30604,g30590,I29204,g31248,g31241,g31257,g27708
	,g31258,g31254,g29966,g31376,g30735,g31514,g31497,g31503
	,g31518,g33066,g32126,g32106,g29195,g31223,g31212,g31228
	,g31188,g30457,g27675,g30459,g31465,g31295,g27880,g32234
	,g32096,g31919,g29952,g27773,g31267,g29043,g27709,g29979
	,I26880,I28567,I28566,g28220,g31931,g27013,g30997,g30999
	,g29982,g29529,g29013,I27314,g31928,g30989,g30996,g30990
	,g31000,I28851,g27998,g31003,g31009,g30337,g30217,g31888
	,g29810,g29789,g29773,g29762,g29743,g29742,g29774,g29693
	,g29799,g31922,g31901,g31913,g27736,g32139,g32113,g33051
	,g29962,g29520,g31885,g31775,I27253,g31911,g31070,g30937
	,g31021,g31554,g31566,g31528,g31672,g31542,g31579,g31710
	,g31170,g31194,g31154,g31327,g30435,g31876,g31908,g30000
	,g32140,g32109,I27232,g27967,g31893,g31468,I27738,g30501
	,I27388,g31904,g30983,g30998,g31770,g31745,g31887,g31918
	,g31773,g31900,g33030,g29311,g29318,g31898,g27774,g30614
	,g30825,g30673,g31912,g33056,I29337,g30309,g29310,g31761
	,g30543,g31316,g31751,g31930,g31881,g31873,g31909,g33020
	,g30305,g30312,g27928,g30522,g27930,g27956,g31781,g33061
	,g27830,g31303,g31279,g31879,g30934,g30929,g31008,g30195
	,g29365,g30578,g30593,g31608,g30572,g31623,g31638,g31653
	,g30567,g33344,g33341,g33364,g33368,g28542,g33340,g33358
	,g33363,g33334,g28228,g33357,g33330,g33333,g33351,g30005
	,g30596,g30592,g28224,g29765,g30568,g30321,g29382,g29755
	,g28231,g29384,g32119,g32145,g29949,g29366,g29373,g31253
	,g31774,g32127,g32107,g30156,g30144,g32017,g31291,g31274
	,g31249,g32108,g30159,g32128,g30148,g32122,g32153,g30150
	,g32103,g30143,g32244,g30130,g31276,g28297,g31767,g32129
	,g32158,g30162,g28141,g30576,g30594,g30589,g30598,g31671
	,g31708,g31326,g30119,g32149,g32159,g30183,g31315,g31308
	,g31269,g32150,g32258,g30302,g30218,g30296,g32151,g32120
	,g30146,g31255,g31320,g32116,g32286,g30171,g31757,g31762
	,g32114,g32146,g30132,g31706,g32104,g30147,g32121,g30134
	,g31306,g31317,g31287,g29147,g31244,g31709,g28336,g28349
	,g31289,g31753,I28832,g28150,g32157,g32143,g30170,g31766
	,g31764,g31768,g31755,g30169,g32148,g32115,g30136,g32147
	,g32248,g30129,g30117,g31284,g31754,g31760,I29013,I29002
	,g30106,g30123,g30160,g28484,g29073,g29192,g28553,g29182
	,g29008,g28528,g28458,I29185,I29182,g28402,g31782,g31785
	,g31749,g28471,g29036,g29188,g28539,g29199,g28982,g29178
	,g29110,g29197,g31325,g29105,g31541,g30157,g32272,g32110
	,g28342,g28659,g28316,g31905,g33025,g28371,I26094,I26367
	,I26050,I26394,I26418,I26460,I26071,I26439,g28357,g31747
	,g28705,g29068,g28497,g28632,g28416,g28404,g29176,g31902
	,g31903,g28698,g31924,g28375,g31889,g28721,g28644,g28707
	,g28731,g28358,g31926,g28435,g28386,g28702,g31914,g28332
	,g32263,g32152,g28295,g28619,g28372,g28286,g28814,g28385
	,g31899,g28618,g28388,g28852,g28750,g31882,g28651,g28305
	,g28335,g30343,g32276,g32112,g32111,g32142,I26419,g31906
	,g28334,g28734,g28691,g31748,g31929,g28629,g28647,g31890
	,g30393,g28646,g31932,g28320,g28728,g31245,g31915,g28348
	,g28649,g28611,g32141,g32156,g31311,g28347,g28640,g28403
	,g31877,g30583,g30573,g30580,g28610,g28665,g28362,g28775
	,g28717,g28609,g28664,I26395,g28361,g31927,g31268,g28662
	,g28685,g28323,g28684,g31923,g31878,g31910,g28635,g31880
	,g30142,g28778,g28727,g31886,g28743,g28428,g28490,g31874
	,g28373,g28329,g31907,g28641,g29938,g31669,g28401,I26461
	,g28328,g28680,g28417,g28344,g28621,g28359,g28600,g31875
	,g28420,g28723,g31302,g28733,g30480,g28390,g28747,g31891
	,g33046,g29166,g28720,g31916,g28815,g28715,g28400,g28776
	,g31892,g28331,g31779,g28816,g33378,g31917,g28308,g28681
	,g30414,g31883,g28306,g31925,g31304,g28716,g28850,g28668
	,g31920,g31921,g31884,g28556,g28530,g33332,g33338,g33342
	,g33327,g33328,g33349,g28239,g33331,g33350,g33355,g33329
	,g33369,g33352,g33372,g33345,g33759,g28249,g33367,g33339
	,g33343,g33362,g28317,g28387,g28628,g28623,g28418,g28682
	,g28744,g28718,g28622,g28345,g28688,g28745,g28310,g28774
	,g28374,g28309,g28319,g31526,I26440,g31259,g28729,g28430
	,g28636,g28772,g28667,g29143,g31260,g28773,g28701,g28296
	,g28746,g28511,g28429,g28719,g28708,g31251,g28749,g28730
	,g28419,g28700,g28732,g28389,g28671,g31772,g28751,g31322
	,g28643,g28634,g32186,g28405,g28851,g28735,g28631,g28322
	,g28704,g28748,g28699,I26072,g28817,g28724,g31473,g28687
	,g28690,g34174,g34084,g31256,g34161,I26368,I26051,g31246
	,g28661,g28650,g28670,g28818,g28884,g28777,I26095,g31466
	,g31250,g33964,g33542,g34071,g33534,g33536,g33539,g33540
	,g34125,g33788,g28588,g33873,g33356,g33361,g34157,g33805
	,g28252,g28571,g33535,g33537,g33732,g33797,g33823,g33717
	,g33710,g33789,g33608,g33733,g30601,g30672,g30237,g30259
	,g30206,g31994,g31989,g31975,g31961,g32302,g32313,g31992
	,g31505,g31944,g32311,g32232,g32281,g32325,g32255,g32290
	,g32008,g32340,g32337,g32270,g32282,I30261,I30192,I29985
	,I30123,I30468,I30054,I30399,I30330,g32118,g32033,g32038
	,g33259,g32030,g33251,g32303,g30609,g32335,g28954,g32328
	,g32410,g32317,I26700,g31933,I26693,g32069,I27481,g32167
	,g31985,g33279,g32013,g32309,g32095,g32161,g32409,g32047
	,g30734,g32266,g32014,g32088,g32056,g33380,g30608,g32082
	,g32054,g31771,g32402,g31941,g30611,I30193,I30055,I29986
	,I30124,g32462,g32534,g32649,g32541,g32613,g32584,g32519
	,g32555,g32476,g32874,g32853,g32713,g32656,g32599,g32504
	,g32548,g32627,g32620,g32881,g32691,g32592,g32634,g32483
	,g32663,g32606,g32684,g32569,g32677,g32469,g32670,g32706
	,g32867,g32527,g32497,g32860,g32888,g32490,g32895,g32562
	,g32902,g32754,g32472,g32573,g32718,g32898,g32927,g32682
	,g32920,g32812,g32833,g32848,g32725,g32515,g32761,g32732
	,g32963,g32653,g32566,g32501,g32588,g32494,g32595,g32617
	,g32559,g32631,g32783,g32458,g32970,g32602,g32696,g32775
	,g32826,g32552,g32710,g32768,g32508,g32949,g32862,g32840
	,g32537,g32891,g32797,g32530,g32905,g32913,g32790,g32703
	,g32523,g32465,g32638,g32747,g32580,g32884,g32487,g32667
	,g32942,g32660,g32624,g32689,g32877,g32819,g32855,g32956
	,g32645,I30400,g32859,g32591,g32612,g32648,g32605,g32683
	,g32554,g32576,g32852,g32518,g32712,g32705,g32489,g32669
	,g32561,g32598,g32887,g32461,g32880,g32533,g32626,g32482
	,g32662,g32583,g32641,g32873,g32475,g32909,g32676,g32468
	,g32619,g32655,g32511,g32866,g32526,g32496,g32894,g32547
	,g32698,g32540,I26682,g32071,g30733,g32097,g32348,g29042
	,g32086,g29372,I26705,g28752,g32342,g32369,g32858,g32946
	,g32788,g32795,g32744,g32758,g32809,g32837,g32939,g32865
	,g32830,g32816,g32823,g32901,g32918,g32967,g32886,g32879
	,g32960,g32737,g32765,g32730,g32802,g32925,g32723,g32932
	,g32872,g32851,g32772,g32751,g32908,g32953,g32633,g32604
	,g32611,g32647,g32640,g32618,g32597,g32590,g32467,g32460
	,g32488,g32474,g32517,g32510,g32503,g32481,g32539,g32525
	,g32532,g32582,g32553,g32575,g32568,g32546,I30331,I30469
	,I30262,g32785,g32777,g32770,g32828,g32972,g32813,g32799
	,g32748,g32915,g32842,g32792,g32958,g32929,g32727,g32806
	,g32720,g32835,g32936,g32922,g32965,g32734,g32763,g32741
	,g32943,g32665,g32693,g32686,g32679,g32672,g32707,g32658
	,g32700,g32628,g32642,g32621,g32635,g32593,g32607,g32614
	,g32600,g32950,g32776,g32719,g32755,g32805,g32798,g32921
	,g32935,g32914,g32733,g32971,g32769,g32827,g32928,g32820
	,g32726,g32834,g32841,g32964,g32762,g32740,g32791,g32784
	,g32957,g32692,g32664,g32678,g32657,g32685,g32714,g32671
	,g32699,g32491,g32463,g32484,g32477,g32470,g32498,g32512
	,g32505,g32563,g32535,g32577,g32570,g32528,g32549,g32542
	,g32556,g32899,g32951,g32849,g32771,g32973,g32906,g32728
	,g32892,g32749,g32836,g32966,g32843,g32856,g32793,g32944
	,g32742,g32786,g32778,g32756,g32821,g32863,g32807,g32814
	,g32800,g32937,g32930,g32721,g32916,g32885,g32923,g32735
	,g32870,g32844,g32871,g32794,g32829,g32729,g32907,g32808
	,g32900,g32864,g32822,g32938,g32893,g32878,g32764,g32736
	,g32924,g32722,g32857,g32959,g32850,g32945,g32779,g32743
	,g32787,g32757,g32750,g32952,g32974,g32815,g32917,g32801
	,g32931,g32473,g32538,g32675,g32567,g32560,g32466,g32704
	,g32524,g32589,g32610,g32668,g32495,g32545,g32459,g32697
	,g32690,g32603,g32646,g32574,g32509,g32711,g32516,g32639
	,g32654,g32531,g32502,g32596,g32480,g32581,g32625,g32661
	,g32632,g33255,g32251,g28779,g32321,g32400,g30605,g30597
	,g32057,I26676,g32414,g33274,I28585,g29539,g32231,g32295
	,I31593,g32099,g32090,I27271,g30591,I28147,g28917,I27784
	,g32200,I26785,g32196,g30317,g28367,I26670,I27777,I26679
	,g32049,I26687,I26649,I28419,g32046,g32191,g32239,g32825
	,g32832,g32767,g32760,g32724,g32789,g32507,g32514,g32500
	,g32962,g32804,g32652,g32934,g32674,g32609,g32883,g32637
	,g32941,g32594,g32630,g32616,g32782,g32623,g32544,g32558
	,g32919,g32955,g32774,g32709,g32869,g32529,g32753,g32681
	,g32811,g32717,g32897,g32890,g32912,g32847,g32904,g32702
	,g32948,g32522,g32464,g32565,g32493,g32746,g32579,g32587
	,g32486,g32479,g32839,g32854,g32876,g32688,g32457,g32695
	,g32818,g32969,g32644,g32659,g32572,g32551,g32739,g32911
	,g32629,g32766,g32701,g32926,g32861,g32521,g32903,g32506
	,g32947,g32940,g32759,g32882,g32745,g32608,g32636,g32622
	,g32485,g32875,g32643,g32954,g32752,g32687,g32571,g32680
	,g32817,g32810,g32471,g32708,g32868,g32499,g32831,g32716
	,g32896,g32961,g32513,g32651,g32803,g32731,g32846,g32933
	,g32673,g32564,g32536,g32796,g32492,g32781,g32615,g32586
	,g32578,g32543,g32478,g32666,g32601,g32557,g32838,g32694
	,g32773,g32550,g32456,g32968,g32824,g32889,g32738,I26664
	,g31596,I27385,g33266,g32224,g30613,g33596,g32188,g33303
	,g30922,g29873,g32198,g30916,g32050,g32356,g31940,g32396
	,g30271,g30315,g30262,g32350,g33597,g33383,g31502,g32310
	,g30252,g33267,g32083,g33254,g32176,g31522,g31943,g33265
	,g33386,g33282,g32067,g33286,g33288,g31189,g33595,g32293
	,g31213,g33277,g33384,g31480,g32376,g32204,g32172,g32072
	,g33272,g33295,g30732,g31495,g32412,g32035,g32203,g33256
	,g33287,g33290,g33297,g32087,g32180,g31496,g32345,I31600
	,g31949,g33271,g32419,g33581,g33298,g33273,g33278,g31959
	,g29730,g30565,g33582,g32250,g30824,g32183,g29725,g29697
	,g33587,I28336,g32084,g32020,g31991,g32265,g32085,g32089
	,g32225,g33393,g32105,g32098,g32018,g31489,g32163,g29286
	,g30458,g32238,I29363,g31273,g31296,g31282,g32170,g32042
	,g32055,g31513,g31871,g33588,g32287,g33598,g31501,g32278
	,g33276,g33590,g31869,g32230,g32070,g33579,g31323,g33270
	,g31283,g31297,g33580,g33589,g29257,g33426,I29149,I27718
	,g30984,I29139,I29368,I27713,g30269,g30284,g30235,g30216
	,g30194,g30226,g32010,g30257,g32009,g29347,g32305,g29326
	,g31967,g30166,g30230,g31986,g30198,g30178,g30188,g30154
	,g32273,g32301,g32306,g29806,g29805,g29842,g29857,g29872
	,g29749,g29766,g29871,g29757,g29783,g29747,g29794,g30001
	,g29758,g32324,g29841,g29856,g29885,g29782,g32323,g32291
	,g30191,g30211,g30190,g30199,g30223,g31968,g31976,g30210
	,g30233,g30272,g30200,g30180,g30243,g31987,g30254,g31237
	,g31242,g31996,g30219,g31966,g31974,g30248,g30208,g30140
	,g30207,g30175,g29320,g30165,g30228,g30152,g30196,g30239
	,g30186,g30185,g31960,g30238,g30229,g30164,g30153,g32269
	,g32330,g32300,g32256,g32241,g29899,g29875,g29874,g29843
	,g32332,g29770,g30024,g32307,g29784,g29807,g29759,g29795
	,g29859,g29751,g29887,g32314,g29785,g32322,g32242,g32292
	,g32312,g30267,g30266,g31993,g30275,g30203,g30234,g30245
	,g29337,g31977,g30246,g30281,g30274,g30192,g31988,g30225
	,g29797,g29798,g32333,g29861,g32326,g29808,g29845,g29909
	,g29788,g29876,g29772,g32315,g29809,g29787,g29891,g32304
	,g29987,g33275,g33387,g33253,g31971,g33268,g29540,g33257
	,g31978,g30282,g29322,g30288,g27925,g30276,g31300,g32175
	,g31286,g31312,g31275,g32171,g31299,g31285,g31950,g33281
	,g29556,g33389,g33390,g29903,g32178,g31321,g31310,g31298
	,g32174,g31309,g31997,g31324,g31314,g32182,g31467,g31301
	,g32179,g31313,g30273,g29315,g30280,g29886,g29316,g29898
	,g30249,g30308,g30260,g33280,g33294,g33292,g29910,g29328
	,g29915,g29900,g29323,g29908,g27380,g31488,g33289,g33293
	,g31266,g32165,g31281,g31272,g27955,g31667,g33296,g27767
	,g30265,g27365,g30240,g32427,g30290,g30316,g30294,g27824
	,g33262,g30285,g33261,g27876,g27401,g29889,g33260,g32408
	,g33571,g31970,g31965,g33604,g33550,g33556,g31942,g31935
	,g29263,g33573,g33606,g29280,g33565,g33572,g33603,g33558
	,g34351,g33605,g33669,g33557,g33548,g33555,g33960,g33250
	,g33574,g33547,g33549,g32398,g29269,g33564,g29292,g30278
	,g30205,g30204,g30289,g30227,g30277,g30268,g30236,g30283
	,g30247,g30258,g30215,g32338,g32283,g32274,g30221,g30250
	,g30231,g30251,g30242,g30241,g30197,g30222,g30209,g30177
	,g30187,g30261,g30167,g32261,g32331,g29750,g29767,g32246
	,g32260,g30264,g30263,g30168,g29331,g30253,g30179,g30244
	,g30232,g30174,g30220,g31990,g29796,g29888,g29760,g29844
	,g29858,g29769,g32343,g32284,g34348,g34146,g30212,g30193
	,g30256,g30255,g30202,g30181,g30224,g30213,g30041,g29860
	,g29890,g29902,g29901,g29771,g29877,g29761,g34322,g34359
	,g34324,g34332,g33566,g29304,g34022,g34069,g34251,g33563
	,g29298,g29222,g33965,g34110,g34111,g33961,g34107,g34147
	,g34073,g34162,g32187,g32194,I29199,g32394,g29041,I29977
	,g32446,g32318,g33134,g33131,g32205,g32990,g28155,g33083
	,I30761,g30182,g33001,g28142,g33000,g32988,g28166,g28162
	,g32994,g29491,g28157,I30734,I28349,g33141,g28262,g33441
	,g29498,I27749,g32999,g33429,g33450,I29582,I30750,g28819
	,I30718,I30746,I30741,I30735,g30328,g31261,g31240,I30728
	,I30756,g28161,g33136,I29913,I30751,g33068,I27735,I31122
	,I31142,I31117,I31087,I31017,I31097,I31032,I31052,I31137
	,I31127,I31042,I31177,I31037,I31082,I31132,I31102,I31162
	,I31167,I31002,I31062,I31027,I31147,I31107,I31092,I31047
	,I31172,I31007,I31072,I31077,I31152,I31057,I31012,I31327
	,I31237,I31317,I31247,I31342,I31202,I31207,I31227,I31197
	,I31337,I31272,I31347,I31277,I31182,I31322,I31192,I31212
	,I31292,I31302,I31332,I31252,I31282,I31307,I31242,I31312
	,I31187,I31257,I31232,I31287,I31297,I31222,I31267,I31352
	,I31262,I31357,I31217,g32520,g32455,I31157,g32585,g32650
	,I31067,I31022,I31112,g32715,g32910,g32780,I27730,g28184
	,I30755,I28838,g33034,I28301,I30727,g33067,g33047,g33060
	,g28163,g32845,I29894,g33054,g31895,g33028,g33052,g32987
	,g32993,I30745,g29185,g28173,g28181,I28540,g33023,g33021
	,g33065,g33385,g33382,g33886,g33863,g33872,g33884,g33857
	,g33866,g33841,g33878,g33943,g33862,g32184,g32189,g32164
	,g32206,g32168,g32177,g32199,g32195,g32193,g33856,g33639
	,g33843,g33877,g33941,g33868,g33837,g33842,g33864,g33855
	,g33869,g33942,g33846,g33860,g33876,g33880,g33887,g33889
	,g33867,g33652,g33861,g29353,g31794,g31479,I29961,g32430
	,g32377,g29358,g31487,I31271,I31316,I31046,I31091,I31136
	,I31001,I31181,I31226,I31296,I31301,I31056,I31016,I31101
	,I31021,I31321,I31071,I31076,I31231,I31326,I31151,I31236
	,I31196,I31261,I31116,I31156,I31121,I31081,I31266,I31201
	,I31341,I31346,I31036,I31306,I31086,I31171,I31041,I31176
	,I31286,I31141,I31311,I31291,I31251,I31006,I31011,I31216
	,I31146,I31061,I31221,I31256,I31066,I31106,I31026,I31111
	,I31241,I31246,I31331,I31031,I31126,I31131,I31336,I31161
	,I31276,I31351,I31166,I31356,I31206,I31281,I31186,I31191
	,I31096,I31211,I31051,g32426,g32357,g31207,g33147,g32353
	,g30914,g33163,g33175,I30717,g33128,g33125,g32347,g31936
	,g33440,g33423,g33312,I29352,g33144,g33139,g33133,g32390
	,g29914,g32352,g32392,I30760,g33138,g33146,g33160,g31969
	,g32388,g31791,g32385,g32387,g33161,g33130,g33135,g30105
	,g33108,I29579,I28866,g32391,g33434,g32336,g32389,g33107
	,g33148,g33145,g33137,g33142,g33100,g32421,I29973,g32442
	,g33143,g33103,g32434,g31945,I29965,g32329,g31218,g31208
	,I30740,g32393,g32359,g33427,g33097,g30411,g33029,g30477
	,g30404,g30399,g33419,g33085,g30398,g33316,g30539,g30397
	,g30441,g30915,g30919,g33009,g33129,g33132,g30465,g30921
	,g30925,g30540,g33048,g30554,g30507,g30412,g33069,g30395
	,g30421,g30430,g33002,g32370,g32986,g30402,g30474,g30413
	,g30401,g32995,g31469,g31373,g30400,g30469,g30434,g30551
	,g30450,g33070,g32362,g32354,g30445,g32346,g30541,g33317
	,g33174,g33162,g33049,g30516,g33447,g33089,g30544,g32997
	,g30511,g32344,g32360,g30462,g33140,g30547,g30531,g32361
	,g32373,g30446,g32991,g30471,g33053,g31231,g31232,g30473
	,g30452,g33062,g30468,g30512,g30447,g30523,g31133,g31127
	,g33055,g30536,g30492,g31372,g31318,g31491,g31483,g33006
	,g32374,I29351,g30518,g30449,g30513,g33304,g33859,g31482
	,g33428,g31476,g33433,g31119,g31117,g31183,g31206,g31220
	,g31224,g33321,g30515,g33432,g33098,g33022,g33315,g33014
	,I29939,g33031,g30563,g33032,g30472,g32349,g32358,g30463
	,g30418,g33057,g33058,g33088,g33093,g32372,g30419,g32996
	,g33449,g33439,g32368,g30410,g31897,g33095,g33096,g30476
	,g33063,g32351,g30396,g30464,g31225,g30533,g30426,g32367
	,g30550,g30467,g30460,g30437,g33017,g30527,g33003,g32386
	,g32992,g30454,g30503,g33024,g32380,g30479,g33033,g30520
	,g30561,g33314,g31498,g31506,g31116,g31068,g32375,g30535
	,g33059,g30491,g33313,g30406,g33437,g32989,g30485,g33094
	,g30425,g30525,g30442,g30422,g30482,g30542,g33010,g30559
	,g30394,g30448,g30508,g30423,g30407,g31507,g32355,g30415
	,g30514,g33018,g30478,g33127,g31896,g32998,g30484,g31229
	,g31226,g30408,g33026,g33084,g30428,g33064,g30433,g30461
	,g30443,g30431,g33050,g31126,g30537,g30500,g30493,g33413
	,g33027,g30417,g30509,g30470,g30409,I28925,g28722,g33849
	,g33647,g28660,g33844,g33640,g33883,g33879,g28327,g33871
	,g33848,g28683,g33106,g28639,g33881,g33865,g33101,g28343
	,g33840,g33858,g28703,g28360,g33882,g33870,g33847,g33885
	,g33646,g33438,g33448,g31121,g33090,g33075,g30926,g33092
	,g34523,g30920,g31515,g32371,g30930,g30927,g33310,g33109
	,g33804,g31219,g31182,g33311,g33305,g31230,g33269,g33264
	,g30495,g33012,g30453,g30496,g30439,g30519,g33007,g30505
	,g30546,g30548,g30403,g30558,g30475,g30429,g30549,g33013
	,g30451,g30488,g33004,g30416,g30545,g34438,g30552,g30517
	,g30529,g30486,g30497,g34524,g34550,g34537,g34048,g30553
	,g30405,g30427,g30489,g30432,g33016,g30560,g30555,g30436
	,g30481,g30502,g30528,g33015,g30534,g30444,g30490,g33005
	,g33011,g30556,g30455,g30510,g30466,g33008,g30562,g30557
	,g30440,g30524,g30521,g30506,g30499,g30532,g30530,g30438
	,g30487,g34543,g30424,g30504,g30526,g30483,g30538,g34252
	,g30494,g32983,g30498,g30420,g34542,g34309,g34330,g34250
	,g34249,g34344,g34346,g34310,g34354,g33039,g31578,g33112
	,g33719,g33237,g33830,g33822,g30295,g33212,g33204,I27567
	,I27576,I28390,g33909,g33910,g32364,g33694,g33487,g33478
	,g33469,g33518,g33515,g33519,g33517,g33516,g33520,g33521
	,g33522,g33523,I27561,g33838,g30072,g30569,I27579,g29368
	,g33197,g33219,g33528,g33506,g33507,g33500,g33502,g33509
	,g33513,g33527,g33512,g33510,g33511,g33524,g33531,g33530
	,g33499,g33503,g33498,g33508,g33525,g33497,g33526,g33504
	,g33501,g33529,g33489,g33493,g33492,g33491,g33490,g33495
	,g33488,g33494,g33484,g33486,g33485,g33479,g33481,g33482
	,g33480,g33496,g33461,g33464,g33463,g33462,g33466,g33468
	,g33467,g33475,g33471,g33477,g33476,g33470,g33473,g33472
	,g29371,g32383,I27549,g33709,g33117,I27742,g32024,g29379
	,I29239,I29236,I27570,g33076,g33381,g30116,I27573,I29245
	,I29248,I27552,I27564,I27555,I28908,I27558,g33326,g32449
	,I27546,g33988,g34018,g33684,g33689,g32117,g33176,g33044
	,g33187,g33685,g33972,g32253,g32267,g33354,g33980,g33976
	,g32437,g33072,g33318,g33979,g33323,g32445,g33430,g34019
	,g33994,g34000,g33149,g33998,g33693,g33700,g34010,g33042
	,g33786,g33706,g33164,g33981,g34011,g34009,g33714,g33703
	,g34017,g34012,g31783,g33969,g33692,g33699,g30606,g32021
	,g33795,g33986,g33041,I28883,g33758,g33968,g33734,g34021
	,I29909,g33676,g33680,g34003,g33036,g33394,g33970,g33532
	,g33505,g33514,g33474,g33465,g33483,g33983,g33040,g33038
	,g33037,g33966,g33043,g33996,g33975,g34002,g34016,g33045
	,g33974,g33967,g33977,g32132,g31591,g33375,g32433,g33421
	,g33412,g33901,g33087,g33722,g33721,g33406,g33411,g33416
	,g33897,g33082,g33405,g33074,g33410,g33401,g33893,g33263
	,g33927,g33718,g33720,g33715,g33408,g33414,g33081,g33896
	,g33404,g33402,g33392,g33446,g33399,g33407,g33073,g33892
	,g33403,g33400,g33418,g33425,g33091,g33904,g33422,g33900
	,g33420,g33086,g33415,g33409,g30991,g33730,g32029,g32031
	,g33832,g33833,g31288,g33911,g33915,g33687,g33681,g32288
	,g32280,g33742,g32032,g32036,g32403,g32411,g33111,g33810
	,g33802,g33690,g33697,g33114,g33809,g33814,g33790,g33787
	,g33760,g32407,g32279,g33784,g32252,g32428,g32420,g33902
	,g33898,g34067,g32294,g33701,g33707,g33785,g32130,g32123
	,g33984,g33811,g33815,g33903,g33905,g32124,g33973,g34005
	,g33995,g29291,g32044,g32045,g33891,g33997,g33908,g33906
	,g32052,g32068,g33982,g32289,g33991,g32039,g32043,g29274
	,g33914,g33835,g33801,g33808,g32240,g32268,g33990,g34015
	,g33834,g33836,g29309,g29262,g33989,g34007,g32048,g32051
	,g29268,g29303,g34004,g32401,g32397,g34014,g32418,g32413
	,g34169,g33541,g33828,g33820,g33922,g33919,g33543,g32131
	,g32144,g34008,g33987,g29297,g29285,g34695,g33993,g34001
	,g33417,g33890,g34702,g34364,g34685,g34698,g34687,g34599
	,g34538,g34535,g34513,g34439,g34545,g34506,g34539,g33807
	,I29891,g33913,g33907,g33616,I30995,g30928,g31666,I28582
	,g34034,I31724,I31727,g31657,I28594,I30641,I30644,g29374
	,I30861,I28591,I31844,I31843,I31838,I31848,I31849,I31854
	,I31853,I31874,I31859,I31873,I31858,I31863,I31864,I31616
	,I31782,I31545,I31459,I31528,I31659,I31770,I31561,I31786
	,I31569,I31486,I31625,I28588,I28872,g34208,g33963,I31869
	,I31868,g34055,g33962,g30155,I31622,I31642,I31482,I31564
	,I31550,I31776,I31539,I31555,I31650,I31779,I31474,I31619
	,I29233,g34082,g34079,g34076,g34083,g33360,g33365,g33239
	,g33796,g34075,g34081,g34078,g34074,g34113,g32028,g31995
	,g33379,I30983,g33431,I29981,g32415,g32450,I30980,g33346
	,g33451,g34148,g34172,g33679,I31839,g33925,g34090,g32381
	,g30729,I30959,I30962,I29936,I29571,I31701,I31686,I31810
	,I31504,I31607,I31800,I31581,g34101,I31610,I31823,I31672
	,I31586,I31807,I31814,I30992,I31817,I31820,I31463,I31466
	,I30986,I31791,I31515,g33686,I31523,g33695,I31597,I31497
	,I31604,I31500,I31803,I31796,I31694,g34099,g33678,g33704
	,g33674,g33728,g33725,g33711,g33675,g33683,g33812,g33819
	,g33831,g33921,g33552,g33575,g33617,g34168,g34006,g34370
	,g33560,g33599,g33578,g33546,g34167,g33545,g33551,g33999
	,g33584,g33586,g33561,g33544,g33992,g34103,g33933,g33930
	,g33585,g34170,g34013,g34231,g33119,g33600,g34026,I30901
	,g33583,g33562,g33607,g34028,g33570,g34193,g33577,g33985
	,g33601,g33553,g33568,g34020,g33554,g33592,g33569,g34100
	,g33602,g33576,g34025,g34190,g33559,g33594,g33116,g33231
	,g33591,g34036,g34035,g33567,g34027,g34095,g34057,g34204
	,g33227,g33978,g32438,g31937,I29969,g33374,g33376,g34117
	,g33242,g33366,g33370,g34226,g34211,g34066,g33359,g33353
	,g33243,g33247,g34774,g33371,g33373,g33249,g33248,g34166
	,g34149,g34158,g34064,g34199,I32352,g33118,g33115,g33238
	,g34206,g34189,g34207,g33234,g33240,g34046,g33236,g34043
	,g34194,g33593,g34440,g34724,g33971,g34742,g34762,g34600
	,g34700,g34693,g34697,g34684,g34703,g34679,g32363,g34024
	,g34291,g31655,g33766,g33641,g33917,g33806,g33708,g33698
	,g33916,g33705,g33713,g33648,g33800,g33772,I28897,g33953
	,g33952,I32364,g30610,g33778,g33653,g33716,g33920,g33712
	,g33912,g33813,g33691,g33631,g33702,g33918,g33761,g33951
	,g33335,I28597,g33080,g32382,g33875,g32384,I29444,g33459
	,g34156,g34181,g34179,g34183,g33620,g33845,g33926,g33929
	,g33665,g33744,g33661,g33736,g33688,g33682,g33621,g34267
	,g33923,g33456,g33637,g33936,g33458,g33934,g33931,g33729
	,g33827,g33937,g33755,g33726,g33928,g33750,g33670,g33932
	,g33839,g33850,g34260,g32015,g32404,g33436,g33609,g34264
	,I29447,g34266,g34261,g34263,I30686,g34268,g33958,g33955
	,g33956,g33954,g34023,g33957,g34262,g34269,g33888,g33454
	,g33424,g32453,g33791,g33455,g33743,g33731,g33803,g34337
	,g34342,g34295,g34341,g34390,g34382,g34385,g34363,g34389
	,g34395,g34410,g34279,g34120,g34173,g34116,g34171,g34394
	,g33798,g34334,g34340,g34338,g33283,g32441,g33442,g33377
	,g34496,g34192,g34132,g34124,g34197,g34053,g34044,g34062
	,g34070,g34068,g34042,g34060,g34049,g33610,g33612,g33618
	,g33624,g34258,g33627,g34257,g33619,g33623,g34790,g33622
	,g33626,g34259,g34345,g33613,g33614,g33625,g33611,g34265
	,g33829,g33818,g34380,g34381,g34365,g34401,g34393,g34281
	,g34414,g34284,g34396,g34415,g34301,g33735,g33821,g33727
	,g33816,g34826,g34842,g34725,g34771,g34741,g34761,g34743
	,g34766,I30766,g34109,g34097,g34102,g34112,g34096,g34087
	,g34086,g34106,g34063,g34212,g34214,g34216,g34213,g34050
	,g34045,g34054,g34230,g34215,g34061,g34104,g34085,g34108
	,g34091,g34065,g34114,g34105,g34186,g34178,g34184,g34182
	,g34180,g34187,g34191,g34185,g33391,g34188,g33388,g33658
	,I31972,I32051,I32109,I31983,I32106,I32062,I29438,g34358
	,g34461,g30917,g34094,I32059,I32119,I32056,I32096,I29585
	,I32158,I32161,g33071,I30998,g33110,g33899,I31829,g33924
	,g34402,g34405,g34319,g33120,g33635,I30971,I32202,I32074
	,I32093,I32079,I32116,g34229,g34047,I32150,g34329,I32185
	,I32067,I32103,I32089,I32071,g34196,g34203,g34205,g34198
	,g34080,g34093,g34072,g34119,g34092,g34115,g34138,g34141
	,g34143,g34217,g34223,g34228,g34225,g34219,g34224,g34218
	,g34098,g34139,g34089,g34088,g34077,g34136,g34133,g34135
	,g34140,g34137,g34253,g34706,g34463,g34465,g34467,g34254
	,g34468,g34037,g34039,g34444,I31535,g34255,g34456,g34462
	,g34449,g34464,g34256,g34443,g34447,g34445,g34446,g34038
	,g34466,g34453,g34029,g34457,I30989,I31491,I31494,g34397
	,g34367,g34388,g34298,g34371,I32639,g34386,g34398,g34335
	,g34287,g34333,g34378,g34375,g34458,g34450,g34441,g34040
	,g34033,g34041,g34448,g34455,g34442,g34032,g34454,g34030
	,g34031,g34452,g34460,g34459,g34451,g34867,g34849,g34791
	,g34819,g34841,g34811,g33228,g34300,g34352,g32027,g34278
	,g34145,g34121,I31973,g34350,g34349,g34160,g34122,I31985
	,I29441,g34321,g34399,g34347,g34314,g34280,g34407,I32607
	,g34353,g34123,g34151,g34152,g34118,I31974,g34282,g34318
	,g34406,g34283,g34412,g34403,g34059,g34416,I31469,g34387
	,I31477,g34404,g34411,g34306,g34305,g34303,g34286,g34323
	,g34326,g34327,g34315,g34313,g34307,g34328,g34336,g34311
	,g34413,g34130,g34142,I32186,g34150,g34126,I32187,I32613
	,g34195,g34275,g34272,g34159,g34134,I32203,g34144,g34131
	,I32204,g33443,g34052,I31361,I32601,I31984,g34153,g33944
	,g33628,g33460,g34202,g34482,g34478,g33660,g33457,g34294
	,g34376,g34331,g34368,g34273,g34274,g33696,g34289,g34372
	,g34421,g34369,g34288,g34293,g34374,g34373,g34290,g34417
	,g34377,g34292,g34379,g34366,g34737,g34297,g34339,g34308
	,g34343,g34312,g34317,g34325,g34320,g34316,g34299,I32651
	,I32654,I32617,I32591,I32621,I32550,I32665,g34569,I32648
	,I32594,I32671,I32645,I32547,g34880,g34866,g34850,g34856
	,I31748,I31751,g34572,g33645,g33638,I32297,g34051,I32222
	,g34420,g34056,g34419,I32231,g34540,I32228,g34271,I32225
	,g34409,I30537,g34558,g34486,g34487,g34479,g34484,g34555
	,g34532,g34556,g34554,g34485,g34476,g34483,g34481,g34529
	,g34527,g34528,g34507,g34509,g34508,g34514,g34526,g34503
	,g34533,g34557,g34534,g34392,I32195,I32192,I32388,I32391
	,g33677,g33657,g34498,g34588,g34582,g34584,g34474,g34536
	,g34580,I32284,g34477,g34475,g34227,I32240,g34408,I32243
	,g34270,g34492,g34494,g34577,I32274,g34544,g34220,I32234
	,g34418,g34400,I32237,g34844,g34497,I31878,g34642,g34637
	,g34058,g34564,g34567,g34568,g34489,g34495,g34493,g34516
	,g34520,g34519,g34525,g34515,g34518,g34517,g34488,g34561
	,g34563,g34566,g34541,g34560,g34562,g34565,g34490,g34499
	,g34573,g34587,g34586,g34470,g34531,g34574,g34571,I32699
	,g34583,g34491,g34553,g34502,g34581,g34578,g34530,g34549
	,g34576,g34585,g34575,g34881,g34909,g33895,g34505,g34242
	,g34522,g34243,I32855,g34244,g34511,I32431,g34512,g34241
	,g34296,I32170,g34708,I32173,g34246,g34501,g34619,g34510
	,g34245,I32439,g34620,g34643,g34627,g34277,g34645,g34636
	,I32788,g34609,g34634,g34624,g34638,g34521,g34248,g34504
	,g34247,I32824,g34641,I32827,g34285,I32794,g34640,g34635
	,g34612,g34633,I32820,g34617,I32803,I32800,g34647,g34644
	,g34646,g34639,g34626,g34611,I32812,g34625,I32837,g34610
	,g34618,g34384,g34222,g34570,g34876,g34686,g34701,g34707
	,g34276,g34127,g34649,g34657,g34630,g34613,g34631,g34602
	,g34621,g34608,g34603,I32806,g34622,g34606,g34601,g34607
	,g34615,g34628,g34614,g34632,g34605,g34598,I32791,I32797
	,I32846,g34616,g34629,g34604,I32782,g34623,I32815,I32809
	,I32843,g34666,g34658,g34662,g34681,g34678,g34661,g34665
	,g34655,g34696,g34710,g34694,g34709,g34911,g34200,g34210
	,I32904,g34209,I32535,I32433,I32452,I32775,I32763,I32461
	,g34699,I32458,I32766,I32455,I32770,g34423,g34559,g34689
	,g34676,g34672,g34673,I32432,g34680,g34670,I32525,g34683
	,g34682,I32440,I32470,I32874,I32473,I32871,g34668,I32476
	,I32464,I32752,I32878,I32467,I32441,g34882,g34732,I32935
	,g34722,I32929,g34719,I32446,I32449,g34715,g34500,g34691
	,g34675,g34677,g34664,g34692,g34671,g34669,g34674,g34720
	,g34726,g34729,g34723,g34721,g34727,g34733,g34735,g34731
	,g34730,g34728,g34734,g34391,g34656,g34428,g34654,g34429
	,I32976,g34430,g34653,g34422,g34659,g34427,g34480,I32305
	,g34736,I32309,g34432,g34716,g34648,g34431,g34424,g34713
	,g34434,g34714,g34433,g34472,g34711,g34471,g34757,g34748
	,g34758,g34763,g34744,g34746,g34756,g34753,g34750,g34426
	,g34755,g34759,g34781,g34745,g34754,g34752,g34765,g34740
	,g34764,g34747,g34751,g34663,I32659,I32516,g34304,I32985
	,g34302,I32840,I32675,I32947,I32960,I32684,g34778,I32681
	,I32956,I32678,I32953,g34667,g34782,I32834,I32693,I32973
	,I32696,I32950,I32687,I32967,I32970,I32690,g34801,g34792
	,g34794,g34803,g34806,g34795,I32991,g34802,g34793,I32988
	,g34805,g34473,I33020,g34799,g34797,g34798,g34804,g34800
	,g34796,g34807,g34808,I32938,g34579,g34769,g34590,g34770
	,g34591,I33053,I33056,g34592,g34772,I32518,g34767,g34589
	,g34690,I32479,g34785,I32482,g34594,g34776,g34775,g34593
	,I32517,g34768,g34596,g34777,g34595,g34688,g34843,g34783
	,g34660,g34786,g34787,g34810,g34760,I32868,g34469,I32884
	,I33027,I33041,g34840,I33037,I33034,I33024,I33075,I32881
	,I33050,I33030,I33044,I33047,I33070,g34738,I32997,g34712
	,g34820,g34823,g34864,g34827,g34813,I32756,g34718,g34833
	,g34830,g34816,g34836,g34717,g34851,g34812,g34848,g34789
	,g34809,I32909,I32757,g34872,g34870,g34868,g34871,g34857
	,g34861,g34859,g34860,g34910,I33067,I33109,I32758,g34862
	,g34863,g34858,g34865,g34874,g34873,g34869,g34875,I33079
	,g34739,I33182,g34650,g34894,g34900,g34890,g34897,g34887
	,g34906,g34884,g34903,g34879,g34847,g34855,I32994,I32921
	,I32963,g34930,I33143,I33146,I33140,I33137,I33134,I33131
	,I33173,I33176,I33155,I33158,I33167,I33170,I33149,I33152
	,I33161,I33164,I33106,I33197,g34773,g34749,g34924,g34920
	,g34926,g34922,g34928,g34914,g34916,g34918,g34878,I32982
	,g34845,g34943,g34934,g34933,g34932,g34942,g34939,g34941
	,g34938,g34940,I33210,g34852,g34784,g34950,g34947,g34951
	,g34949,g34952,g34944,g34945,g34946,I33064,I33119,g34883
	,g34954,g34967,g34964,g34961,g34966,g34968,g34962,g34965
	,g34963,g34912,I33214,g34893,g34846,g34977,g34970,g34975
	,g34978,g34979,g34971,g34976,g34974,I33103,I33179,g34931
	,I33264,I33255,I33246,I33261,I33252,I33258,I33249,I33267
	,g34929,g34877,g34955,g34987,g34982,g34985,g34988,g34989
	,g34983,g34986,g34984,I33189,I33285,I33276,I33270,I33282
	,I33218,I33273,I33279,I33291,I33288,g34935,g34960,g34994
	,g34990,g34992,g34995,g34996,g34997,g34993,g34991,g34953
	,g34948,g34969,g34957,g34980,I33235,I33232,g34973,g34981
	,g34998,g34999,g35000,I33297,g35001,I33300,g35002;

	dff 	XG1 	(g5057,g33046);
	dff 	XG2 	(g2771,g34441);
	dff 	XG3 	(g1882,g33982);
	dff 	XG4 	(g6462,g25751);
	dff 	XG5 	(g2299,g34007);
	dff 	XG6 	(g4040,g24276);
	dff 	XG7 	(g2547,g30381);
	dff 	XG8 	(g559,g640);
	dff 	XG9 	(g640,g637);
	dff 	XG10 	(g3017,g31877);
	dff 	XG11 	(g3243,g30405);
	dff 	XG12 	(g452,g25604);
	dff 	XG13 	(g464,g25607);
	dff 	XG14 	(g3542,g30416);
	dff 	XG15 	(g5232,g30466);
	dff 	XG16 	(g5813,g25736);
	dff 	XG17 	(g2907,g34617);
	dff 	XG18 	(g1744,g33974);
	dff 	XG19 	(g5909,g30505);
	dff 	XG20 	(g1802,g33554);
	dff 	XG21 	(g3554,g30432);
	dff 	XG22 	(g6219,g33064);
	dff 	XG23 	(g807,g34881);
	dff 	XG24 	(g6031,g6027);
	dff 	XG25 	(g6027,g6023);
	dff 	XG26 	(g847,g24216);
	dff 	XG27 	(g976,g24232);
	dff 	XG28 	(g4172,g34733);
	dff 	XG29 	(g4372,g34882);
	dff 	XG30 	(g3512,g33026);
	dff 	XG31 	(g749,g31867);
	dff 	XG32 	(g3490,g25668);
	dff 	XG33 	(g6005,g24344);
	dff 	XG34 	(g4235,g4232);
	dff 	XG35 	(g4232,g4229);
	dff 	XG36 	(g1600,g33966);
	dff 	XG37 	(g1714,g33550);
	dff 	XG38 	(g3649,g3625);
	dff 	XG39 	(g3625,g3618);
	dff 	XG40 	(g3155,g30393);
	dff 	XG41 	(g3355,g31880);
	dff 	XG42 	(g2236,g29248);
	dff 	XG43 	(g4555,g4571);
	dff 	XG44 	(g4571,g6974);
	dff 	XG45 	(g3698,g24274);
	dff 	XG46 	(g6073,g31920);
	dff 	XG47 	(g1736,g33973);
	dff 	XG48 	(g1968,g30360);
	dff 	XG49 	(g4621,g34460);
	dff 	XG50 	(g5607,g30494);
	dff 	XG51 	(g2657,g30384);
	dff 	XG52 	(g5659,g24340);
	dff 	XG53 	(g490,g29223);
	dff 	XG54 	(g311,g26881);
	dff 	XG55 	(g6069,g31925);
	dff 	XG56 	(g772,g34252);
	dff 	XG57 	(g5587,g30489);
	dff 	XG58 	(g6177,g29301);
	dff 	XG59 	(g6377,g6373);
	dff 	XG60 	(g6373,g6369);
	dff 	XG61 	(g3167,g33022);
	dff 	XG62 	(g5615,g30496);
	dff 	XG63 	(g4567,g33043);
	dff 	XG64 	(g3057,g28062);
	dff 	XG65 	(g3457,g29263);
	dff 	XG66 	(g6287,g30533);
	dff 	XG67 	(g1500,g24256);
	dff 	XG68 	(g2563,g34015);
	dff 	XG69 	(g4776,g34031);
	dff 	XG70 	(g4593,g34452);
	dff 	XG71 	(g6199,g34646);
	dff 	XG72 	(g2295,g34001);
	dff 	XG73 	(g1384,g25633);
	dff 	XG74 	(g1339,g24259);
	dff 	XG75 	(g5180,g33049);
	dff 	XG76 	(g2844,g34609);
	dff 	XG77 	(g1024,g31869);
	dff 	XG78 	(g5591,g30490);
	dff 	XG79 	(g3598,g30427);
	dff 	XG80 	(g4264,g21894);
	dff 	XG81 	(g767,g33965);
	dff 	XG82 	(g5853,g34645);
	dff 	XG83 	(g3321,g3317);
	dff 	XG84 	(g3317,g3298);
	dff 	XG85 	(g2089,g33571);
	dff 	XG86 	(g4933,g34267);
	dff 	XG87 	(g4521,g26971);
	dff 	XG88 	(g5507,g34644);
	dff 	XG89 	(g3618,g3661);
	dff 	XG90 	(g6291,g30534);
	dff 	XG91 	(g294,g33535);
	dff 	XG92 	(g5559,g30498);
	dff 	XG93 	(g5794,g25728);
	dff 	XG94 	(g6144,g25743);
	dff 	XG95 	(g3813,g25684);
	dff 	XG96 	(g562,g25613);
	dff 	XG97 	(g608,g34438);
	dff 	XG98 	(g1205,g24244);
	dff 	XG99 	(g3909,g30439);
	dff 	XG100 	(g6259,g30541);
	dff 	XG101 	(g5905,g30519);
	dff 	XG102 	(g921,g25621);
	dff 	XG103 	(g2955,g34807);
	dff 	XG104 	(g203,g25599);
	dff 	XG105 	(g6088,g31924);
	dff 	XG106 	(g1099,g24235);
	dff 	XG107 	(g4878,g34036);
	dff 	XG108 	(g5204,g30476);
	dff 	XG109 	(g5630,g5623);
	dff 	XG110 	(g5623,g5666);
	dff 	XG111 	(g3606,g30429);
	dff 	XG112 	(g1926,g32997);
	dff 	XG113 	(g6215,g33063);
	dff 	XG114 	(g3586,g30424);
	dff 	XG115 	(g291,g32977);
	dff 	XG116 	(g4674,g34026);
	dff 	XG117 	(g3570,g30420);
	dff 	XG118 	(g637,g24212);
	dff 	XG119 	(g5969,g6012);
	dff 	XG120 	(g6012,g5983);
	dff 	XG121 	(g1862,g33560);
	dff 	XG122 	(g676,g29226);
	dff 	XG123 	(g843,g25619);
	dff 	XG124 	(g4132,g28076);
	dff 	XG125 	(g4332,g34455);
	dff 	XG126 	(g4153,g30457);
	dff 	XG127 	(g5666,g5637);
	dff 	XG128 	(g5637,g5659);
	dff 	XG129 	(g6336,g33625);
	dff 	XG130 	(g622,g34790);
	dff 	XG131 	(g3506,g30414);
	dff 	XG132 	(g4558,g26966);
	dff 	XG133 	(g6065,g31923);
	dff 	XG134 	(g6322,g6315);
	dff 	XG135 	(g6315,g6358);
	dff 	XG136 	(g3111,g25656);
	dff 	XG137 	(g117,g30390);
	dff 	XG138 	(g2837,g26935);
	dff 	XG139 	(g939,g34727);
	dff 	XG140 	(g278,g25594);
	dff 	XG141 	(g4492,g26963);
	dff 	XG142 	(g4864,g34034);
	dff 	XG143 	(g1036,g33541);
	dff 	XG144 	(g128,g28093);
	dff 	XG145 	(g1178,g24236);
	dff 	XG146 	(g3239,g30404);
	dff 	XG147 	(g718,g28051);
	dff 	XG148 	(g6195,g29303);
	dff 	XG149 	(g1135,g26917);
	dff 	XG150 	(g6137,g25741);
	dff 	XG151 	(g6395,g33624);
	dff 	XG152 	(g3380,g31882);
	dff 	XG153 	(g5343,g24337);
	dff 	XG154 	(g554,g34911);
	dff 	XG155 	(g496,g33963);
	dff 	XG156 	(g3853,g34627);
	dff 	XG157 	(g5134,g29282);
	dff 	XG158 	(g1422,g1418);
	dff 	XG159 	(g1418,g24254);
	dff 	XG160 	(g3794,g25676);
	dff 	XG161 	(g2485,g33013);
	dff 	XG162 	(g925,g32981);
	dff 	XG163 	(g48,g34993);
	dff 	XG164 	(g5555,g30483);
	dff 	XG165 	(g878,g875);
	dff 	XG166 	(g875,g869);
	dff 	XG167 	(g1798,g32994);
	dff 	XG168 	(g4076,g28070);
	dff 	XG169 	(g2941,g34806);
	dff 	XG170 	(g3905,g30453);
	dff 	XG171 	(g763,g33539);
	dff 	XG172 	(g6255,g30526);
	dff 	XG173 	(g4375,g26951);
	dff 	XG174 	(g4871,g34035);
	dff 	XG175 	(g4722,g34636);
	dff 	XG176 	(g590,g32978);
	dff 	XG177 	(g6692,g6668);
	dff 	XG178 	(g6668,g6661);
	dff 	XG179 	(g1632,g30348);
	dff 	XG180 	(g5313,g24336);
	dff 	XG181 	(g3100,g3092);
	dff 	XG182 	(g3092,g25648);
	dff 	XG183 	(g1495,g24250);
	dff 	XG184 	(g6497,g6490);
	dff 	XG185 	(g6490,g25757);
	dff 	XG186 	(g1437,g29236);
	dff 	XG187 	(g6154,g29298);
	dff 	XG188 	(g1579,g1576);
	dff 	XG189 	(g1576,g24255);
	dff 	XG190 	(g5567,g30499);
	dff 	XG191 	(g1752,g33976);
	dff 	XG192 	(g1917,g32996);
	dff 	XG193 	(g744,g30335);
	dff 	XG194 	(g3040,g31878);
	dff 	XG195 	(g4737,g34637);
	dff 	XG196 	(g4809,g25693);
	dff 	XG197 	(g6267,g30528);
	dff 	XG198 	(g3440,g25661);
	dff 	XG199 	(g3969,g4012);
	dff 	XG200 	(g4012,g3983);
	dff 	XG201 	(g1442,g24251);
	dff 	XG202 	(g5965,g30521);
	dff 	XG203 	(g4477,g26960);
	dff 	XG204 	(g1233,g24239);
	dff 	XG205 	(g4643,g34259);
	dff 	XG206 	(g5264,g30474);
	dff 	XG207 	(g6329,g6351);
	dff 	XG208 	(g6351,g24348);
	dff 	XG209 	(g2610,g33016);
	dff 	XG210 	(g5160,g34643);
	dff 	XG211 	(g5360,g31905);
	dff 	XG212 	(g5933,g30510);
	dff 	XG213 	(g1454,g29239);
	dff 	XG214 	(g753,g26897);
	dff 	XG215 	(g1296,g34729);
	dff 	XG216 	(g3151,g34625);
	dff 	XG217 	(g2980,g34800);
	dff 	XG218 	(g6727,g24353);
	dff 	XG219 	(g3530,g33029);
	dff 	XG220 	(g4742,g21903);
	dff 	XG221 	(g4104,g33615);
	dff 	XG222 	(g1532,g24253);
	dff 	XG223 	(g4304,g24281);
	dff 	XG224 	(g2177,g33997);
	dff 	XG225 	(g3010,g25651);
	dff 	XG226 	(g52,g34997);
	dff 	XG227 	(g4754,g34263);
	dff 	XG228 	(g1189,g24237);
	dff 	XG229 	(g2287,g33584);
	dff 	XG230 	(g4273,g24280);
	dff 	XG231 	(g1389,g26920);
	dff 	XG232 	(g1706,g33548);
	dff 	XG233 	(g5835,g29296);
	dff 	XG234 	(g1171,g30338);
	dff 	XG235 	(g4269,g21895);
	dff 	XG236 	(g2399,g33588);
	dff 	XG237 	(g3372,g31886);
	dff 	XG238 	(g4983,g34041);
	dff 	XG239 	(g5611,g30495);
	dff 	XG240 	(g3661,g3632);
	dff 	XG241 	(g4572,g29279);
	dff 	XG242 	(g3143,g25655);
	dff 	XG243 	(g2898,g34795);
	dff 	XG244 	(g3343,g24269);
	dff 	XG245 	(g3235,g30403);
	dff 	XG246 	(g4543,g33042);
	dff 	XG247 	(g3566,g30419);
	dff 	XG248 	(g4534,g34023);
	dff 	XG249 	(g4961,g28090);
	dff 	XG250 	(g6398,g31926);
	dff 	XG251 	(g4927,g34642);
	dff 	XG252 	(g2259,g30370);
	dff 	XG253 	(g2819,g34448);
	dff 	XG254 	(g4414,g26946);
	dff 	XG255 	(g5802,g5794);
	dff 	XG256 	(g2852,g34610);
	dff 	XG257 	(g417,g24209);
	dff 	XG258 	(g681,g28047);
	dff 	XG259 	(g437,g24206);
	dff 	XG260 	(g351,g26891);
	dff 	XG261 	(g5901,g30504);
	dff 	XG262 	(g2886,g34798);
	dff 	XG263 	(g3494,g25669);
	dff 	XG264 	(g5511,g30480);
	dff 	XG265 	(g3518,g33027);
	dff 	XG266 	(g1604,g33972);
	dff 	XG267 	(g4135,g28077);
	dff 	XG268 	(g5092,g25697);
	dff 	XG269 	(g4831,g28099);
	dff 	XG270 	(g4382,g26947);
	dff 	XG271 	(g6386,g24350);
	dff 	XG272 	(g479,g24210);
	dff 	XG273 	(g3965,g30455);
	dff 	XG274 	(g4749,g28084);
	dff 	XG275 	(g2008,g33993);
	dff 	XG276 	(g736,g802);
	dff 	XG277 	(g802,g799);
	dff 	XG278 	(g3933,g30444);
	dff 	XG279 	(g222,g33537);
	dff 	XG280 	(g3050,g25650);
	dff 	XG281 	(g5736,g31915);
	dff 	XG282 	(g1052,g25625);
	dff 	XG283 	(g58,g30328);
	dff 	XG284 	(g2122,g30366);
	dff 	XG285 	(g2465,g33593);
	dff 	XG286 	(g6483,g25755);
	dff 	XG287 	(g5889,g30502);
	dff 	XG288 	(g4495,g33036);
	dff 	XG289 	(g365,g25595);
	dff 	XG290 	(g4653,g34462);
	dff 	XG291 	(g3179,g33024);
	dff 	XG292 	(g1728,g33552);
	dff 	XG293 	(g2433,g34014);
	dff 	XG294 	(g3835,g29273);
	dff 	XG295 	(g6187,g25748);
	dff 	XG296 	(g4917,g34638);
	dff 	XG297 	(g1070,g30341);
	dff 	XG298 	(g822,g26899);
	dff 	XG299 	(g6023,g6019);
	dff 	XG300 	(g914,g30336);
	dff 	XG301 	(g5339,g5335);
	dff 	XG302 	(g5335,g5331);
	dff 	XG303 	(g4164,g26940);
	dff 	XG304 	(g969,g25622);
	dff 	XG305 	(g2807,g34447);
	dff 	XG306 	(g5424,g25709);
	dff 	XG307 	(g4054,g33613);
	dff 	XG308 	(g6191,g25749);
	dff 	XG309 	(g5077,g25704);
	dff 	XG310 	(g5523,g33053);
	dff 	XG311 	(g3680,g3676);
	dff 	XG312 	(g3676,g3672);
	dff 	XG313 	(g6637,g30555);
	dff 	XG314 	(g174,g25601);
	dff 	XG315 	(g1682,g33971);
	dff 	XG316 	(g355,g26892);
	dff 	XG317 	(g1087,g1083);
	dff 	XG318 	(g1083,g1079);
	dff 	XG319 	(g1105,g26915);
	dff 	XG320 	(g2342,g33008);
	dff 	XG321 	(g6307,g30538);
	dff 	XG322 	(g3802,g3794);
	dff 	XG323 	(g6159,g25750);
	dff 	XG324 	(g2255,g30369);
	dff 	XG325 	(g2815,g34446);
	dff 	XG326 	(g911,g29230);
	dff 	XG327 	(g43,g34789);
	dff 	XG328 	(g3983,g4005);
	dff 	XG329 	(g1748,g33975);
	dff 	XG330 	(g5551,g30497);
	dff 	XG331 	(g5742,g31917);
	dff 	XG332 	(g3558,g30418);
	dff 	XG333 	(g5499,g25721);
	dff 	XG334 	(g2960,g34622);
	dff 	XG335 	(g3901,g30438);
	dff 	XG336 	(g4888,g34266);
	dff 	XG337 	(g6251,g30540);
	dff 	XG338 	(g6358,g6329);
	dff 	XG339 	(g1373,g32986);
	dff 	XG340 	(g157,g33960);
	dff 	XG341 	(g2783,g34442);
	dff 	XG342 	(g4281,g4277);
	dff 	XG343 	(g4277,g21896);
	dff 	XG344 	(g3574,g30421);
	dff 	XG345 	(g2112,g33573);
	dff 	XG346 	(g1283,g34730);
	dff 	XG347 	(g433,g24205);
	dff 	XG348 	(g4297,g4294);
	dff 	XG349 	(g4294,g21900);
	dff 	XG350 	(g5983,g6005);
	dff 	XG351 	(g1459,g1399);
	dff 	XG352 	(g1399,g24257);
	dff 	XG353 	(g758,g32979);
	dff 	XG354 	(g5712,g25731);
	dff 	XG355 	(g4138,g28078);
	dff 	XG356 	(g4639,g34025);
	dff 	XG357 	(g6537,g25763);
	dff 	XG358 	(g5543,g30481);
	dff 	XG359 	(g1582,g1500);
	dff 	XG360 	(g3736,g31890);
	dff 	XG361 	(g5961,g30517);
	dff 	XG362 	(g6243,g30539);
	dff 	XG363 	(g632,g34880);
	dff 	XG364 	(g1227,g24242);
	dff 	XG365 	(g3889,g30436);
	dff 	XG366 	(g3476,g29265);
	dff 	XG367 	(g1664,g32990);
	dff 	XG368 	(g1246,g24245);
	dff 	XG369 	(g6128,g25739);
	dff 	XG370 	(g6629,g30553);
	dff 	XG371 	(g246,g26907);
	dff 	XG372 	(g4049,g24278);
	dff 	XG373 	(g4449,g26955);
	dff 	XG374 	(g2932,g24282);
	dff 	XG375 	(g4575,g29276);
	dff 	XG376 	(g4098,g31894);
	dff 	XG377 	(g4498,g33037);
	dff 	XG378 	(g528,g26894);
	dff 	XG379 	(g5436,g25711);
	dff 	XG380 	(g16,g34593);
	dff 	XG381 	(g3139,g25654);
	dff 	XG382 	(g102,g33962);
	dff 	XG383 	(g4584,g34451);
	dff 	XG384 	(g142,g34250);
	dff 	XG385 	(g5331,g5327);
	dff 	XG386 	(g5831,g29295);
	dff 	XG387 	(g239,g26905);
	dff 	XG388 	(g1216,g25629);
	dff 	XG389 	(g2848,g34792);
	dff 	XG390 	(g5805,g5798);
	dff 	XG391 	(g5798,g25729);
	dff 	XG392 	(g5022,g25703);
	dff 	XG393 	(g4019,g4000);
	dff 	XG394 	(g4000,g3976);
	dff 	XG395 	(g1030,g32983);
	dff 	XG396 	(g3672,g3668);
	dff 	XG397 	(g3668,g3649);
	dff 	XG398 	(g3231,g30402);
	dff 	XG399 	(g1430,g1426);
	dff 	XG400 	(g1426,g1422);
	dff 	XG401 	(g4452,g4446);
	dff 	XG402 	(g4446,g26954);
	dff 	XG403 	(g2241,g33999);
	dff 	XG404 	(g1564,g24262);
	dff 	XG405 	(g6148,g6140);
	dff 	XG406 	(g6140,g25742);
	dff 	XG407 	(g6649,g30558);
	dff 	XG408 	(g110,g34848);
	dff 	XG409 	(g884,g881);
	dff 	XG410 	(g881,g878);
	dff 	XG411 	(g3742,g31892);
	dff 	XG412 	(g225,g26901);
	dff 	XG413 	(g4486,g26961);
	dff 	XG414 	(g4504,g33039);
	dff 	XG415 	(g5873,g33059);
	dff 	XG416 	(g5037,g31899);
	dff 	XG417 	(g2319,g33007);
	dff 	XG418 	(g5495,g25720);
	dff 	XG419 	(g4185,g21891);
	dff 	XG420 	(g5208,g30462);
	dff 	XG421 	(g2152,g18422);
	dff 	XG422 	(g5579,g30487);
	dff 	XG423 	(g5869,g33058);
	dff 	XG424 	(g5719,g31916);
	dff 	XG425 	(g1589,g24261);
	dff 	XG426 	(g5752,g25730);
	dff 	XG427 	(g6279,g30531);
	dff 	XG428 	(g5917,g30506);
	dff 	XG429 	(g2975,g34804);
	dff 	XG430 	(g6167,g25747);
	dff 	XG431 	(g4005,g24275);
	dff 	XG432 	(g2599,g33601);
	dff 	XG433 	(g1448,g26922);
	dff 	XG434 	(g3712,g25679);
	dff 	XG435 	(g2370,g29250);
	dff 	XG436 	(g5164,g30459);
	dff 	XG437 	(g1333,g1582);
	dff 	XG438 	(g153,g33534);
	dff 	XG439 	(g6549,g30543);
	dff 	XG440 	(g4087,g29275);
	dff 	XG441 	(g4801,g34030);
	dff 	XG442 	(g2984,g34980);
	dff 	XG443 	(g3961,g30451);
	dff 	XG444 	(g5770,g25723);
	dff 	XG445 	(g962,g25627);
	dff 	XG446 	(g101,g34787);
	dff 	XG447 	(g4226,g4222);
	dff 	XG448 	(g4222,g4219);
	dff 	XG449 	(g6625,g30552);
	dff 	XG450 	(g51,g34996);
	dff 	XG451 	(g1018,g30337);
	dff 	XG452 	(g4045,g24277);
	dff 	XG453 	(g1467,g29237);
	dff 	XG454 	(g2461,g30378);
	dff 	XG455 	(g5706,g31912);
	dff 	XG456 	(g457,g25603);
	dff 	XG457 	(g2756,g33019);
	dff 	XG458 	(g5990,g33623);
	dff 	XG459 	(g471,g25608);
	dff 	XG460 	(g1256,g29235);
	dff 	XG461 	(g5029,g31902);
	dff 	XG462 	(g6519,g29306);
	dff 	XG463 	(g4169,g28080);
	dff 	XG464 	(g1816,g33978);
	dff 	XG465 	(g4369,g26970);
	dff 	XG466 	(g3436,g25660);
	dff 	XG467 	(g5787,g25726);
	dff 	XG468 	(g4578,g29278);
	dff 	XG469 	(g4459,g34253);
	dff 	XG470 	(g3831,g29272);
	dff 	XG471 	(g2514,g33595);
	dff 	XG472 	(g3288,g33610);
	dff 	XG473 	(g2403,g33589);
	dff 	XG474 	(g2145,g34605);
	dff 	XG475 	(g1700,g30350);
	dff 	XG476 	(g513,g25611);
	dff 	XG477 	(g2841,g26936);
	dff 	XG478 	(g5297,g33619);
	dff 	XG479 	(g3805,g3798);
	dff 	XG480 	(g3798,g25677);
	dff 	XG481 	(g2763,g34022);
	dff 	XG482 	(g4793,g34033);
	dff 	XG483 	(g952,g34726);
	dff 	XG484 	(g1263,g31870);
	dff 	XG485 	(g1950,g33985);
	dff 	XG486 	(g5138,g29283);
	dff 	XG487 	(g2307,g34003);
	dff 	XG488 	(g5109,g5101);
	dff 	XG489 	(g5101,g25700);
	dff 	XG490 	(g5791,g25727);
	dff 	XG491 	(g4664,g34463);
	dff 	XG492 	(g2223,g33006);
	dff 	XG493 	(g5808,g29292);
	dff 	XG494 	(g6645,g30557);
	dff 	XG495 	(g2016,g33989);
	dff 	XG496 	(g5759,g28098);
	dff 	XG497 	(g3873,g33033);
	dff 	XG498 	(g3632,g3654);
	dff 	XG499 	(g3654,g24271);
	dff 	XG500 	(g2315,g34005);
	dff 	XG501 	(g2811,g26932);
	dff 	XG502 	(g5957,g30516);
	dff 	XG503 	(g2047,g33575);
	dff 	XG504 	(g3869,g33032);
	dff 	XG505 	(g3719,g31891);
	dff 	XG506 	(g5575,g30486);
	dff 	XG507 	(g46,g34991);
	dff 	XG508 	(g3752,g25678);
	dff 	XG509 	(g3917,g30440);
	dff 	XG510 	(g4188,g4191);
	dff 	XG511 	(g4191,g21901);
	dff 	XG512 	(g1585,g1570);
	dff 	XG513 	(g1570,g24258);
	dff 	XG514 	(g4388,g26949);
	dff 	XG515 	(g6275,g30530);
	dff 	XG516 	(g6311,g30542);
	dff 	XG517 	(g4216,g4213);
	dff 	XG518 	(g4213,g4185);
	dff 	XG519 	(g1041,g25624);
	dff 	XG520 	(g2595,g30383);
	dff 	XG521 	(g2537,g33597);
	dff 	XG522 	(g136,g34598);
	dff 	XG523 	(g4430,g26957);
	dff 	XG524 	(g4564,g26967);
	dff 	XG525 	(g3454,g3447);
	dff 	XG526 	(g3447,g25663);
	dff 	XG527 	(g4826,g28102);
	dff 	XG528 	(g6239,g30524);
	dff 	XG529 	(g3770,g25671);
	dff 	XG530 	(g232,g26903);
	dff 	XG531 	(g5268,g30475);
	dff 	XG532 	(g6545,g34647);
	dff 	XG533 	(g2417,g30377);
	dff 	XG534 	(g1772,g33553);
	dff 	XG535 	(g4741,g21902);
	dff 	XG536 	(g5052,g31903);
	dff 	XG537 	(g5452,g25715);
	dff 	XG538 	(g1890,g33984);
	dff 	XG539 	(g2629,g33602);
	dff 	XG540 	(g572,g28045);
	dff 	XG541 	(g2130,g34603);
	dff 	XG542 	(g4108,g33035);
	dff 	XG543 	(g4308,g4304);
	dff 	XG544 	(g475,g24208);
	dff 	XG545 	(g990,g1239);
	dff 	XG546 	(g1239,g1157);
	dff 	XG547 	(g31,g34596);
	dff 	XG548 	(g3412,g28064);
	dff 	XG549 	(g45,g34990);
	dff 	XG550 	(g799,g24213);
	dff 	XG551 	(g3706,g31887);
	dff 	XG552 	(g3990,g33614);
	dff 	XG553 	(g5385,g31907);
	dff 	XG554 	(g5881,g33060);
	dff 	XG555 	(g1992,g30362);
	dff 	XG556 	(g3029,g31875);
	dff 	XG557 	(g3171,g33023);
	dff 	XG558 	(g3787,g25674);
	dff 	XG559 	(g812,g26898);
	dff 	XG560 	(g832,g25618);
	dff 	XG561 	(g5897,g30518);
	dff 	XG562 	(g4165,g28079);
	dff 	XG563 	(g3281,g3303);
	dff 	XG564 	(g3303,g24267);
	dff 	XG565 	(g4455,g26959);
	dff 	XG566 	(g2902,g34801);
	dff 	XG567 	(g333,g26884);
	dff 	XG568 	(g168,g25600);
	dff 	XG569 	(g2823,g26933);
	dff 	XG570 	(g3684,g28066);
	dff 	XG571 	(g3639,g33612);
	dff 	XG572 	(g5327,g5308);
	dff 	XG573 	(g3338,g24268);
	dff 	XG574 	(g5406,g25716);
	dff 	XG575 	(g3791,g25675);
	dff 	XG576 	(g269,g26906);
	dff 	XG577 	(g401,g24203);
	dff 	XG578 	(g6040,g24346);
	dff 	XG579 	(g441,g24207);
	dff 	XG580 	(g5105,g25701);
	dff 	XG581 	(g3808,g29269);
	dff 	XG582 	(g9,g34592);
	dff 	XG583 	(g3759,g28068);
	dff 	XG584 	(g4467,g34255);
	dff 	XG585 	(g3957,g30450);
	dff 	XG586 	(g4093,g30456);
	dff 	XG587 	(g1760,g32991);
	dff 	XG588 	(g6151,g6144);
	dff 	XG589 	(g160,g34249);
	dff 	XG590 	(g5445,g25713);
	dff 	XG591 	(g5373,g31909);
	dff 	XG592 	(g2279,g30371);
	dff 	XG593 	(g3498,g29268);
	dff 	XG594 	(g586,g29224);
	dff 	XG595 	(g869,g859);
	dff 	XG596 	(g859,g26900);
	dff 	XG597 	(g2619,g33017);
	dff 	XG598 	(g1183,g30339);
	dff 	XG599 	(g1608,g33967);
	dff 	XG600 	(g4197,g4194);
	dff 	XG601 	(g4194,g4188);
	dff 	XG602 	(g5283,g5276);
	dff 	XG603 	(g5276,g5320);
	dff 	XG604 	(g1779,g33559);
	dff 	XG605 	(g2652,g29255);
	dff 	XG606 	(g5459,g5452);
	dff 	XG607 	(g2193,g30368);
	dff 	XG608 	(g2393,g30375);
	dff 	XG609 	(g5767,g25732);
	dff 	XG610 	(g661,g28052);
	dff 	XG611 	(g4950,g28089);
	dff 	XG612 	(g5535,g33055);
	dff 	XG613 	(g2834,g30392);
	dff 	XG614 	(g1361,g30343);
	dff 	XG615 	(g3419,g25657);
	dff 	XG616 	(g6235,g30523);
	dff 	XG617 	(g1146,g24233);
	dff 	XG618 	(g2625,g33018);
	dff 	XG619 	(g150,g32976);
	dff 	XG620 	(g1696,g30349);
	dff 	XG621 	(g6555,g33067);
	dff 	XG622 	(g3385,g31883);
	dff 	XG623 	(g3881,g33034);
	dff 	XG624 	(g6621,g30551);
	dff 	XG625 	(g3470,g25667);
	dff 	XG626 	(g3897,g30452);
	dff 	XG627 	(g518,g25612);
	dff 	XG628 	(g3025,g31874);
	dff 	XG629 	(g538,g34719);
	dff 	XG630 	(g2606,g33607);
	dff 	XG631 	(g1472,g26923);
	dff 	XG632 	(g6113,g25746);
	dff 	XG633 	(g542,g24211);
	dff 	XG634 	(g5188,g33050);
	dff 	XG635 	(g5689,g24341);
	dff 	XG636 	(g1116,g1056);
	dff 	XG637 	(g1056,g24241);
	dff 	XG638 	(g405,g24201);
	dff 	XG639 	(g5216,g30463);
	dff 	XG640 	(g6494,g6486);
	dff 	XG641 	(g6486,g25756);
	dff 	XG642 	(g4669,g34464);
	dff 	XG643 	(g5428,g25710);
	dff 	XG644 	(g996,g24243);
	dff 	XG645 	(g4531,g24335);
	dff 	XG646 	(g2860,g34611);
	dff 	XG647 	(g4743,g34262);
	dff 	XG648 	(g6593,g30546);
	dff 	XG649 	(g2710,g18527);
	dff 	XG650 	(g215,g25591);
	dff 	XG651 	(g4411,g4414);
	dff 	XG652 	(g1413,g30347);
	dff 	XG653 	(g4474,g10384);
	dff 	XG654 	(g5308,g5283);
	dff 	XG655 	(g6641,g30556);
	dff 	XG656 	(g3045,g33020);
	dff 	XG657 	(g6,g34589);
	dff 	XG658 	(g1936,g33562);
	dff 	XG659 	(g55,g35002);
	dff 	XG660 	(g504,g25610);
	dff 	XG661 	(g2587,g33015);
	dff 	XG662 	(g4480,g31896);
	dff 	XG663 	(g2311,g34004);
	dff 	XG664 	(g3602,g30428);
	dff 	XG665 	(g5571,g30485);
	dff 	XG666 	(g3578,g30422);
	dff 	XG667 	(g468,g25606);
	dff 	XG668 	(g5448,g25714);
	dff 	XG669 	(g3767,g25680);
	dff 	XG670 	(g5827,g29294);
	dff 	XG671 	(g3582,g30423);
	dff 	XG672 	(g6271,g30529);
	dff 	XG673 	(g4688,g34028);
	dff 	XG674 	(g5774,g25724);
	dff 	XG675 	(g2380,g33587);
	dff 	XG676 	(g5196,g30460);
	dff 	XG677 	(g5396,g31910);
	dff 	XG678 	(g3227,g30401);
	dff 	XG679 	(g2020,g33990);
	dff 	XG680 	(g3976,g3969);
	dff 	XG681 	(g1079,g1075);
	dff 	XG682 	(g1075,g24238);
	dff 	XG683 	(g6541,g29309);
	dff 	XG684 	(g3203,g30411);
	dff 	XG685 	(g1668,g33546);
	dff 	XG686 	(g4760,g28085);
	dff 	XG687 	(g262,g26904);
	dff 	XG688 	(g1840,g33556);
	dff 	XG689 	(g70,g18093);
	dff 	XG690 	(g5467,g25722);
	dff 	XG691 	(g460,g25605);
	dff 	XG692 	(g6209,g33062);
	dff 	XG693 	(g74,g26893);
	dff 	XG694 	(g5290,g5313);
	dff 	XG695 	(g655,g28050);
	dff 	XG696 	(g3502,g34626);
	dff 	XG697 	(g2204,g33583);
	dff 	XG698 	(g5256,g30472);
	dff 	XG699 	(g4608,g34454);
	dff 	XG700 	(g794,g34850);
	dff 	XG701 	(g4023,g4019);
	dff 	XG702 	(g4423,g4537);
	dff 	XG703 	(g4537,g34024);
	dff 	XG704 	(g3689,g24272);
	dff 	XG705 	(g5381,g31906);
	dff 	XG706 	(g5685,g5681);
	dff 	XG707 	(g5681,g5677);
	dff 	XG708 	(g703,g24214);
	dff 	XG709 	(g5421,g25718);
	dff 	XG710 	(g862,g26909);
	dff 	XG711 	(g3247,g30406);
	dff 	XG712 	(g2040,g33569);
	dff 	XG713 	(g4999,g25694);
	dff 	XG714 	(g4146,g34628);
	dff 	XG715 	(g4633,g34458);
	dff 	XG716 	(g1157,g24240);
	dff 	XG717 	(g5723,g31918);
	dff 	XG718 	(g4732,g34634);
	dff 	XG719 	(g5817,g29293);
	dff 	XG720 	(g2151,g18421);
	dff 	XG721 	(g2351,g33009);
	dff 	XG722 	(g2648,g33603);
	dff 	XG723 	(g6736,g24355);
	dff 	XG724 	(g4944,g34268);
	dff 	XG725 	(g4072,g25691);
	dff 	XG726 	(g344,g26890);
	dff 	XG727 	(g4443,g4449);
	dff 	XG728 	(g3466,g29264);
	dff 	XG729 	(g4116,g28072);
	dff 	XG730 	(g5041,g31900);
	dff 	XG731 	(g5441,g25712);
	dff 	XG732 	(g4434,g26956);
	dff 	XG733 	(g3827,g29271);
	dff 	XG734 	(g6500,g29304);
	dff 	XG735 	(g5673,g5654);
	dff 	XG736 	(g5654,g5630);
	dff 	XG737 	(g3133,g29261);
	dff 	XG738 	(g3333,g28063);
	dff 	XG739 	(g979,g1116);
	dff 	XG740 	(g4681,g34027);
	dff 	XG741 	(g298,g33961);
	dff 	XG742 	(g3774,g25672);
	dff 	XG743 	(g2667,g33604);
	dff 	XG744 	(g3396,g33025);
	dff 	XG745 	(g4210,g4207);
	dff 	XG746 	(g4207,g4204);
	dff 	XG747 	(g1894,g32995);
	dff 	XG748 	(g2988,g34624);
	dff 	XG749 	(g3538,g30415);
	dff 	XG750 	(g301,g33536);
	dff 	XG751 	(g341,g26888);
	dff 	XG752 	(g827,g28055);
	dff 	XG753 	(g6077,g31921);
	dff 	XG754 	(g2555,g33600);
	dff 	XG755 	(g5011,g28105);
	dff 	XG756 	(g199,g34721);
	dff 	XG757 	(g6523,g29307);
	dff 	XG758 	(g1526,g30345);
	dff 	XG759 	(g4601,g34453);
	dff 	XG760 	(g854,g32980);
	dff 	XG761 	(g1484,g29238);
	dff 	XG762 	(g4922,g34639);
	dff 	XG763 	(g5080,g25695);
	dff 	XG764 	(g5863,g33057);
	dff 	XG765 	(g4581,g26969);
	dff 	XG766 	(g3021,g31879);
	dff 	XG767 	(g2518,g29253);
	dff 	XG768 	(g2567,g34021);
	dff 	XG769 	(g568,g26895);
	dff 	XG770 	(g3263,g30413);
	dff 	XG771 	(g6613,g30549);
	dff 	XG772 	(g6044,g24347);
	dff 	XG773 	(g6444,g25758);
	dff 	XG774 	(g2965,g34808);
	dff 	XG775 	(g5857,g30501);
	dff 	XG776 	(g1616,g33969);
	dff 	XG777 	(g890,g34440);
	dff 	XG778 	(g5976,g5969);
	dff 	XG779 	(g3562,g30433);
	dff 	XG780 	(g1404,g26921);
	dff 	XG781 	(g3723,g31893);
	dff 	XG782 	(g3817,g29270);
	dff 	XG783 	(g93,g34878);
	dff 	XG784 	(g4501,g33038);
	dff 	XG785 	(g287,g31865);
	dff 	XG786 	(g2724,g26926);
	dff 	XG787 	(g4704,g28083);
	dff 	XG788 	(g22,g29209);
	dff 	XG789 	(g2878,g34797);
	dff 	XG790 	(g5220,g30478);
	dff 	XG791 	(g617,g34724);
	dff 	XG792 	(g316,g26883);
	dff 	XG793 	(g1277,g32985);
	dff 	XG794 	(g6513,g25761);
	dff 	XG795 	(g336,g26886);
	dff 	XG796 	(g2882,g34796);
	dff 	XG797 	(g933,g32982);
	dff 	XG798 	(g1906,g33561);
	dff 	XG799 	(g305,g26880);
	dff 	XG800 	(g8,g34591);
	dff 	XG801 	(g3368,g31884);
	dff 	XG802 	(g2799,g26931);
	dff 	XG803 	(g887,g884);
	dff 	XG804 	(g4912,g34641);
	dff 	XG805 	(g4157,g34629);
	dff 	XG806 	(g2541,g33598);
	dff 	XG807 	(g2153,g33576);
	dff 	XG808 	(g550,g34720);
	dff 	XG809 	(g255,g26902);
	dff 	XG810 	(g1945,g29244);
	dff 	XG811 	(g5240,g30468);
	dff 	XG812 	(g1478,g26924);
	dff 	XG813 	(g3080,g25645);
	dff 	XG814 	(g3863,g33031);
	dff 	XG815 	(g1959,g29245);
	dff 	XG816 	(g3480,g29266);
	dff 	XG817 	(g6653,g30559);
	dff 	XG818 	(g6719,g6715);
	dff 	XG819 	(g6715,g6711);
	dff 	XG820 	(g2864,g34794);
	dff 	XG821 	(g4894,g28087);
	dff 	XG822 	(g5677,g5673);
	dff 	XG823 	(g3857,g30435);
	dff 	XG824 	(g499,g25609);
	dff 	XG825 	(g5413,g28095);
	dff 	XG826 	(g1002,g28057);
	dff 	XG827 	(g776,g34439);
	dff 	XG828 	(g28,g34595);
	dff 	XG829 	(g1236,g1233);
	dff 	XG830 	(g4646,g34260);
	dff 	XG831 	(g2476,g33012);
	dff 	XG832 	(g1657,g32989);
	dff 	XG833 	(g2375,g34006);
	dff 	XG834 	(g63,g34847);
	dff 	XG835 	(g358,g365);
	dff 	XG836 	(g896,g26910);
	dff 	XG837 	(g967,g21722);
	dff 	XG838 	(g3423,g25658);
	dff 	XG839 	(g283,g28043);
	dff 	XG840 	(g3161,g33021);
	dff 	XG841 	(g2384,g29251);
	dff 	XG842 	(g3361,g25665);
	dff 	XG843 	(g6675,g6697);
	dff 	XG844 	(g6697,g24352);
	dff 	XG845 	(g4616,g34456);
	dff 	XG846 	(g4561,g26968);
	dff 	XG847 	(g2024,g33991);
	dff 	XG848 	(g3451,g3443);
	dff 	XG849 	(g3443,g25662);
	dff 	XG850 	(g2795,g26930);
	dff 	XG851 	(g613,g34599);
	dff 	XG852 	(g4527,g28082);
	dff 	XG853 	(g1844,g33557);
	dff 	XG854 	(g5937,g30511);
	dff 	XG855 	(g4546,g33045);
	dff 	XG856 	(g3103,g3096);
	dff 	XG857 	(g3096,g25649);
	dff 	XG858 	(g2523,g30379);
	dff 	XG859 	(g2643,g34020);
	dff 	XG860 	(g6109,g28100);
	dff 	XG861 	(g1489,g24249);
	dff 	XG862 	(g5390,g31908);
	dff 	XG863 	(g194,g25592);
	dff 	XG864 	(g2551,g30382);
	dff 	XG865 	(g5156,g29285);
	dff 	XG866 	(g3072,g25644);
	dff 	XG867 	(g1242,g1227);
	dff 	XG868 	(g47,g34992);
	dff 	XG869 	(g1955,g33563);
	dff 	XG870 	(g6049,g33622);
	dff 	XG871 	(g3034,g31876);
	dff 	XG872 	(g2273,g33582);
	dff 	XG873 	(g6711,g6692);
	dff 	XG874 	(g4771,g28086);
	dff 	XG875 	(g6098,g25744);
	dff 	XG876 	(g3147,g29262);
	dff 	XG877 	(g3347,g24270);
	dff 	XG878 	(g2269,g33581);
	dff 	XG879 	(g191,g194);
	dff 	XG880 	(g2712,g26937);
	dff 	XG881 	(g626,g34849);
	dff 	XG882 	(g2729,g28060);
	dff 	XG883 	(g5357,g33618);
	dff 	XG884 	(g4991,g34038);
	dff 	XG885 	(g6019,g6000);
	dff 	XG886 	(g6000,g5976);
	dff 	XG887 	(g4709,g34032);
	dff 	XG888 	(g6419,g31927);
	dff 	XG889 	(g6052,g31919);
	dff 	XG890 	(g2927,g34803);
	dff 	XG891 	(g4340,g34459);
	dff 	XG892 	(g5929,g30509);
	dff 	XG893 	(g4907,g34640);
	dff 	XG894 	(g3298,g3274);
	dff 	XG895 	(g4035,g28069);
	dff 	XG896 	(g2946,g21899);
	dff 	XG897 	(g918,g31868);
	dff 	XG898 	(g4082,g26938);
	dff 	XG899 	(g2036,g30363);
	dff 	XG900 	(g577,g30334);
	dff 	XG901 	(g1620,g33970);
	dff 	XG902 	(g2831,g30391);
	dff 	XG903 	(g667,g25615);
	dff 	XG904 	(g930,g33540);
	dff 	XG905 	(g3937,g30445);
	dff 	XG906 	(g5782,g25725);
	dff 	XG907 	(g817,g25617);
	dff 	XG908 	(g1249,g24247);
	dff 	XG909 	(g837,g24215);
	dff 	XG910 	(g599,g33964);
	dff 	XG911 	(g5475,g25719);
	dff 	XG912 	(g739,g29228);
	dff 	XG913 	(g5949,g30514);
	dff 	XG914 	(g6682,g33627);
	dff 	XG915 	(g6105,g28101);
	dff 	XG916 	(g904,g24231);
	dff 	XG917 	(g2873,g34615);
	dff 	XG918 	(g1854,g30356);
	dff 	XG919 	(g5084,g25696);
	dff 	XG920 	(g5603,g30493);
	dff 	XG921 	(g4219,g4216);
	dff 	XG922 	(g2495,g33594);
	dff 	XG923 	(g2437,g34009);
	dff 	XG924 	(g2102,g30365);
	dff 	XG925 	(g2208,g33004);
	dff 	XG926 	(g2579,g34018);
	dff 	XG927 	(g4064,g25685);
	dff 	XG928 	(g4899,g34040);
	dff 	XG929 	(g2719,g25639);
	dff 	XG930 	(g4785,g34029);
	dff 	XG931 	(g5583,g30488);
	dff 	XG932 	(g781,g34600);
	dff 	XG933 	(g6173,g29300);
	dff 	XG934 	(g6369,g6365);
	dff 	XG935 	(g2917,g34802);
	dff 	XG936 	(g686,g25614);
	dff 	XG937 	(g1252,g28058);
	dff 	XG938 	(g671,g29225);
	dff 	XG939 	(g2265,g33580);
	dff 	XG940 	(g6283,g30532);
	dff 	XG941 	(g6365,g6346);
	dff 	XG942 	(g5320,g5290);
	dff 	XG943 	(g6459,g25760);
	dff 	XG944 	(g901,g25620);
	dff 	XG945 	(g5527,g33054);
	dff 	XG946 	(g4489,g26962);
	dff 	XG947 	(g1974,g33564);
	dff 	XG948 	(g1270,g32984);
	dff 	XG949 	(g4966,g34039);
	dff 	XG950 	(g6415,g31932);
	dff 	XG951 	(g6227,g33065);
	dff 	XG952 	(g3929,g30443);
	dff 	XG953 	(g5503,g29291);
	dff 	XG954 	(g4242,g24279);
	dff 	XG955 	(g5925,g30508);
	dff 	XG956 	(g1124,g29232);
	dff 	XG957 	(g4955,g34269);
	dff 	XG958 	(g5224,g30464);
	dff 	XG959 	(g2012,g33988);
	dff 	XG960 	(g6203,g30522);
	dff 	XG961 	(g5120,g25708);
	dff 	XG962 	(g2389,g30374);
	dff 	XG963 	(g4438,g26953);
	dff 	XG964 	(g2429,g34008);
	dff 	XG965 	(g2787,g34444);
	dff 	XG966 	(g1287,g34731);
	dff 	XG967 	(g2675,g33606);
	dff 	XG968 	(g66,g24334);
	dff 	XG969 	(g4836,g34265);
	dff 	XG970 	(g1199,g30340);
	dff 	XG971 	(g5547,g30482);
	dff 	XG972 	(g3782,g25673);
	dff 	XG973 	(g6428,g31929);
	dff 	XG974 	(g2138,g34604);
	dff 	XG975 	(g2338,g33591);
	dff 	XG976 	(g4229,g4226);
	dff 	XG977 	(g6247,g30525);
	dff 	XG978 	(g2791,g26929);
	dff 	XG979 	(g3949,g30448);
	dff 	XG980 	(g1291,g34602);
	dff 	XG981 	(g5945,g30513);
	dff 	XG982 	(g5244,g30469);
	dff 	XG983 	(g2759,g33608);
	dff 	XG984 	(g6741,g33626);
	dff 	XG985 	(g785,g34725);
	dff 	XG986 	(g1259,g30342);
	dff 	XG987 	(g3484,g29267);
	dff 	XG988 	(g209,g25593);
	dff 	XG989 	(g6609,g30548);
	dff 	XG990 	(g5517,g33052);
	dff 	XG991 	(g2449,g34012);
	dff 	XG992 	(g2575,g34017);
	dff 	XG993 	(g65,g34785);
	dff 	XG994 	(g2715,g24263);
	dff 	XG995 	(g936,g26912);
	dff 	XG996 	(g2098,g30364);
	dff 	XG997 	(g4462,g34254);
	dff 	XG998 	(g604,g34251);
	dff 	XG999 	(g6589,g30560);
	dff 	XG1000 	(g1886,g33983);
	dff 	XG1001 	(g6466,g25752);
	dff 	XG1002 	(g6346,g6322);
	dff 	XG1003 	(g429,g24204);
	dff 	XG1004 	(g1870,g33980);
	dff 	XG1005 	(g4249,g34631);
	dff 	XG1006 	(g6455,g28103);
	dff 	XG1007 	(g3004,g31873);
	dff 	XG1008 	(g1825,g29243);
	dff 	XG1009 	(g6133,g25740);
	dff 	XG1010 	(g1008,g25623);
	dff 	XG1011 	(g4392,g26950);
	dff 	XG1012 	(g5002,g4999);
	dff 	XG1013 	(g3546,g30431);
	dff 	XG1014 	(g5236,g30467);
	dff 	XG1015 	(g1768,g30353);
	dff 	XG1016 	(g4854,g34467);
	dff 	XG1017 	(g3925,g30442);
	dff 	XG1018 	(g6509,g29305);
	dff 	XG1019 	(g732,g25616);
	dff 	XG1020 	(g2504,g29252);
	dff 	XG1021 	(g1322,g1459);
	dff 	XG1022 	(g4520,g6972);
	dff 	XG1023 	(g2185,g33003);
	dff 	XG1024 	(g37,g34613);
	dff 	XG1025 	(g4031,g4027);
	dff 	XG1026 	(g4027,g4023);
	dff 	XG1027 	(g2070,g33570);
	dff 	XG1028 	(g4812,g4809);
	dff 	XG1029 	(g6093,g33061);
	dff 	XG1030 	(g968,g21723);
	dff 	XG1031 	(g4176,g34734);
	dff 	XG1032 	(g4405,g4408);
	dff 	XG1033 	(g4408,g26945);
	dff 	XG1034 	(g872,g887);
	dff 	XG1035 	(g6181,g29302);
	dff 	XG1036 	(g6381,g24349);
	dff 	XG1037 	(g4765,g34264);
	dff 	XG1038 	(g5563,g30484);
	dff 	XG1039 	(g1395,g25634);
	dff 	XG1040 	(g1913,g33567);
	dff 	XG1041 	(g2331,g33585);
	dff 	XG1042 	(g6263,g30527);
	dff 	XG1043 	(g50,g34995);
	dff 	XG1044 	(g3945,g30447);
	dff 	XG1045 	(g347,g344);
	dff 	XG1046 	(g5731,g31914);
	dff 	XG1047 	(g4473,g34256);
	dff 	XG1048 	(g1266,g25630);
	dff 	XG1049 	(g5489,g29290);
	dff 	XG1050 	(g714,g29227);
	dff 	XG1051 	(g2748,g31872);
	dff 	XG1052 	(g5471,g29287);
	dff 	XG1053 	(g4540,g31897);
	dff 	XG1054 	(g6723,g6719);
	dff 	XG1055 	(g6605,g30562);
	dff 	XG1056 	(g2445,g34011);
	dff 	XG1057 	(g2173,g33996);
	dff 	XG1058 	(g4287,g21898);
	dff 	XG1059 	(g2491,g33014);
	dff 	XG1060 	(g4849,g34465);
	dff 	XG1061 	(g2169,g33995);
	dff 	XG1062 	(g2283,g30372);
	dff 	XG1063 	(g6585,g30545);
	dff 	XG1064 	(g121,g30389);
	dff 	XG1065 	(g2407,g33590);
	dff 	XG1066 	(g2868,g34616);
	dff 	XG1067 	(g2767,g26927);
	dff 	XG1068 	(g1783,g32992);
	dff 	XG1069 	(g3310,g3281);
	dff 	XG1070 	(g1312,g25631);
	dff 	XG1071 	(g5212,g30477);
	dff 	XG1072 	(g4245,g34632);
	dff 	XG1073 	(g645,g28046);
	dff 	XG1074 	(g4291,g4287);
	dff 	XG1075 	(g79,g26896);
	dff 	XG1076 	(g182,g25602);
	dff 	XG1077 	(g1129,g26916);
	dff 	XG1078 	(g2227,g33578);
	dff 	XG1079 	(g6058,g25745);
	dff 	XG1080 	(g4204,g4200);
	dff 	XG1081 	(g2246,g33579);
	dff 	XG1082 	(g1830,g30354);
	dff 	XG1083 	(g3590,g30425);
	dff 	XG1084 	(g392,g24200);
	dff 	XG1085 	(g1592,g33544);
	dff 	XG1086 	(g6505,g25764);
	dff 	XG1087 	(g6411,g31930);
	dff 	XG1088 	(g1221,g24246);
	dff 	XG1089 	(g5921,g30507);
	dff 	XG1090 	(g106,g26889);
	dff 	XG1091 	(g146,g30333);
	dff 	XG1092 	(g218,g215);
	dff 	XG1093 	(g6474,g25753);
	dff 	XG1094 	(g1932,g32998);
	dff 	XG1095 	(g1624,g32987);
	dff 	XG1096 	(g5062,g25702);
	dff 	XG1097 	(g5462,g29286);
	dff 	XG1098 	(g2689,g34606);
	dff 	XG1099 	(g6573,g33070);
	dff 	XG1100 	(g1677,g29240);
	dff 	XG1101 	(g2028,g32999);
	dff 	XG1102 	(g2671,g33605);
	dff 	XG1103 	(g34,g34877);
	dff 	XG1104 	(g1848,g33558);
	dff 	XG1105 	(g3089,g25647);
	dff 	XG1106 	(g3731,g31889);
	dff 	XG1107 	(g86,g25699);
	dff 	XG1108 	(g5485,g29289);
	dff 	XG1109 	(g2741,g30388);
	dff 	XG1110 	(g2638,g29254);
	dff 	XG1111 	(g4122,g28074);
	dff 	XG1112 	(g4322,g34450);
	dff 	XG1113 	(g5941,g30512);
	dff 	XG1114 	(g2108,g33572);
	dff 	XG1115 	(g25,g15048);
	dff 	XG1116 	(g1644,g33551);
	dff 	XG1117 	(g595,g33538);
	dff 	XG1118 	(g2217,g33005);
	dff 	XG1119 	(g1319,g24248);
	dff 	XG1120 	(g2066,g33002);
	dff 	XG1121 	(g1152,g24234);
	dff 	XG1122 	(g5252,g30471);
	dff 	XG1123 	(g2165,g34000);
	dff 	XG1124 	(g2571,g34016);
	dff 	XG1125 	(g5176,g33048);
	dff 	XG1126 	(g391,g26911);
	dff 	XG1127 	(g5005,g5002);
	dff 	XG1128 	(g2711,g18528);
	dff 	XG1129 	(g1211,g25628);
	dff 	XG1130 	(g2827,g26934);
	dff 	XG1131 	(g6423,g31928);
	dff 	XG1132 	(g4859,g34468);
	dff 	XG1133 	(g424,g24202);
	dff 	XG1134 	(g1274,g33542);
	dff 	XG1135 	(g85,g34717);
	dff 	XG1136 	(g2803,g34445);
	dff 	XG1137 	(g6451,g28104);
	dff 	XG1138 	(g1821,g33555);
	dff 	XG1139 	(g2509,g34013);
	dff 	XG1140 	(g5073,g28091);
	dff 	XG1141 	(g1280,g26919);
	dff 	XG1142 	(g4815,g4812);
	dff 	XG1143 	(g6633,g30554);
	dff 	XG1144 	(g5124,g29281);
	dff 	XG1145 	(g6303,g30537);
	dff 	XG1146 	(g5069,g28092);
	dff 	XG1147 	(g2994,g34732);
	dff 	XG1148 	(g650,g28049);
	dff 	XG1149 	(g1636,g33545);
	dff 	XG1150 	(g3921,g30441);
	dff 	XG1151 	(g2093,g29247);
	dff 	XG1152 	(g6732,g24354);
	dff 	XG1153 	(g1306,g25636);
	dff 	XG1154 	(g5377,g31911);
	dff 	XG1155 	(g1061,g26914);
	dff 	XG1156 	(g3462,g25670);
	dff 	XG1157 	(g2181,g33998);
	dff 	XG1158 	(g956,g25626);
	dff 	XG1159 	(g1756,g33977);
	dff 	XG1160 	(g5849,g29297);
	dff 	XG1161 	(g4112,g28071);
	dff 	XG1162 	(g2685,g30387);
	dff 	XG1163 	(g2197,g33577);
	dff 	XG1164 	(g6116,g25737);
	dff 	XG1165 	(g2421,g33592);
	dff 	XG1166 	(g1046,g26913);
	dff 	XG1167 	(g482,g28044);
	dff 	XG1168 	(g4401,g26948);
	dff 	XG1169 	(g6434,g31931);
	dff 	XG1170 	(g1514,g30344);
	dff 	XG1171 	(g329,g26885);
	dff 	XG1172 	(g6565,g33069);
	dff 	XG1173 	(g2950,g34621);
	dff 	XG1174 	(g4129,g28075);
	dff 	XG1175 	(g1345,g28059);
	dff 	XG1176 	(g6533,g25762);
	dff 	XG1177 	(g3274,g3267);
	dff 	XG1178 	(g3085,g25646);
	dff 	XG1179 	(g4727,g34633);
	dff 	XG1180 	(g1536,g26925);
	dff 	XG1181 	(g3941,g30446);
	dff 	XG1182 	(g370,g25597);
	dff 	XG1183 	(g5694,g24342);
	dff 	XG1184 	(g1858,g30357);
	dff 	XG1185 	(g446,g26908);
	dff 	XG1186 	(g4932,g21905);
	dff 	XG1187 	(g3219,g30399);
	dff 	XG1188 	(g1811,g29242);
	dff 	XG1189 	(g3431,g25659);
	dff 	XG1190 	(g6601,g30547);
	dff 	XG1191 	(g3376,g31881);
	dff 	XG1192 	(g2441,g34010);
	dff 	XG1193 	(g1874,g33986);
	dff 	XG1194 	(g4349,g34257);
	dff 	XG1195 	(g6581,g30544);
	dff 	XG1196 	(g6597,g30561);
	dff 	XG1197 	(g5008,g5005);
	dff 	XG1198 	(g3610,g30430);
	dff 	XG1199 	(g2890,g34799);
	dff 	XG1200 	(g1978,g33565);
	dff 	XG1201 	(g1612,g33968);
	dff 	XG1202 	(g112,g34879);
	dff 	XG1203 	(g2856,g34793);
	dff 	XG1204 	(g6479,g25754);
	dff 	XG1205 	(g1982,g33566);
	dff 	XG1206 	(g6661,g6704);
	dff 	XG1207 	(g5228,g30465);
	dff 	XG1208 	(g4119,g28073);
	dff 	XG1209 	(g6390,g24351);
	dff 	XG1210 	(g1542,g30346);
	dff 	XG1211 	(g4258,g21893);
	dff 	XG1212 	(g4818,g4815);
	dff 	XG1213 	(g5033,g31904);
	dff 	XG1214 	(g4717,g34635);
	dff 	XG1215 	(g1554,g25637);
	dff 	XG1216 	(g3849,g29274);
	dff 	XG1217 	(g6704,g6675);
	dff 	XG1218 	(g3199,g30396);
	dff 	XG1219 	(g5845,g25735);
	dff 	XG1220 	(g4975,g34037);
	dff 	XG1221 	(g790,g34791);
	dff 	XG1222 	(g5913,g30520);
	dff 	XG1223 	(g1902,g30358);
	dff 	XG1224 	(g6163,g29299);
	dff 	XG1225 	(g4125,g28081);
	dff 	XG1226 	(g4821,g28096);
	dff 	XG1227 	(g4939,g28088);
	dff 	XG1228 	(g3207,g30397);
	dff 	XG1229 	(g4483,g4520);
	dff 	XG1230 	(g3259,g30409);
	dff 	XG1231 	(g5142,g29284);
	dff 	XG1232 	(g5248,g30470);
	dff 	XG1233 	(g2126,g30367);
	dff 	XG1234 	(g3694,g24273);
	dff 	XG1235 	(g5481,g29288);
	dff 	XG1236 	(g1964,g30359);
	dff 	XG1237 	(g5097,g25698);
	dff 	XG1238 	(g3215,g30398);
	dff 	XG1239 	(g111,g34718);
	dff 	XG1240 	(g4427,g26952);
	dff 	XG1241 	(g7,g34590);
	dff 	XG1242 	(g2779,g26928);
	dff 	XG1243 	(g4200,g4197);
	dff 	XG1244 	(g1720,g30351);
	dff 	XG1245 	(g1367,g31871);
	dff 	XG1246 	(g5112,g5105);
	dff 	XG1247 	(g19,g34594);
	dff 	XG1248 	(g4145,g26939);
	dff 	XG1249 	(g2161,g33994);
	dff 	XG1250 	(g376,g25596);
	dff 	XG1251 	(g2361,g33586);
	dff 	XG1252 	(g582,g31866);
	dff 	XG1253 	(g2051,g33000);
	dff 	XG1254 	(g1193,g26918);
	dff 	XG1255 	(g5401,g33051);
	dff 	XG1256 	(g3408,g28065);
	dff 	XG1257 	(g2327,g30373);
	dff 	XG1258 	(g907,g28056);
	dff 	XG1259 	(g947,g34601);
	dff 	XG1260 	(g1834,g30355);
	dff 	XG1261 	(g3594,g30426);
	dff 	XG1262 	(g2999,g34805);
	dff 	XG1263 	(g5727,g31913);
	dff 	XG1264 	(g2303,g34002);
	dff 	XG1265 	(g3065,g25652);
	dff 	XG1266 	(g699,g28053);
	dff 	XG1267 	(g723,g29229);
	dff 	XG1268 	(g5703,g33620);
	dff 	XG1269 	(g546,g34722);
	dff 	XG1270 	(g2472,g33599);
	dff 	XG1271 	(g5953,g30515);
	dff 	XG1272 	(g6439,g33066);
	dff 	XG1273 	(g1740,g33979);
	dff 	XG1274 	(g3550,g30417);
	dff 	XG1275 	(g3845,g25683);
	dff 	XG1276 	(g2116,g33574);
	dff 	XG1277 	(g3195,g30410);
	dff 	XG1278 	(g3913,g30454);
	dff 	XG1279 	(g1687,g33547);
	dff 	XG1280 	(g2681,g30386);
	dff 	XG1281 	(g2533,g33596);
	dff 	XG1282 	(g324,g26887);
	dff 	XG1283 	(g2697,g34607);
	dff 	XG1284 	(g5747,g33056);
	dff 	XG1285 	(g4417,g31895);
	dff 	XG1286 	(g6561,g33068);
	dff 	XG1287 	(g1141,g29233);
	dff 	XG1288 	(g2413,g30376);
	dff 	XG1289 	(g1710,g33549);
	dff 	XG1290 	(g6527,g29308);
	dff 	XG1291 	(g6404,g25759);
	dff 	XG1292 	(g3255,g30408);
	dff 	XG1293 	(g1691,g29241);
	dff 	XG1294 	(g2936,g34620);
	dff 	XG1295 	(g5644,g33621);
	dff 	XG1296 	(g5152,g25707);
	dff 	XG1297 	(g5352,g24339);
	dff 	XG1298 	(g6120,g25738);
	dff 	XG1299 	(g2775,g34443);
	dff 	XG1300 	(g2922,g34619);
	dff 	XG1301 	(g1111,g29234);
	dff 	XG1302 	(g5893,g30503);
	dff 	XG1303 	(g1311,g21724);
	dff 	XG1304 	(g3267,g3310);
	dff 	XG1305 	(g6617,g30550);
	dff 	XG1306 	(g2060,g33001);
	dff 	XG1307 	(g4512,g33040);
	dff 	XG1308 	(g5599,g30492);
	dff 	XG1309 	(g3401,g25664);
	dff 	XG1310 	(g4366,g26944);
	dff 	XG1311 	(g94,g34614);
	dff 	XG1312 	(g3129,g29260);
	dff 	XG1313 	(g3329,g3325);
	dff 	XG1314 	(g3325,g3321);
	dff 	XG1315 	(g5170,g33047);
	dff 	XG1316 	(g4456,g25692);
	dff 	XG1317 	(g5821,g25733);
	dff 	XG1318 	(g6299,g30536);
	dff 	XG1319 	(g3727,g31888);
	dff 	XG1320 	(g2079,g29246);
	dff 	XG1321 	(g4698,g34261);
	dff 	XG1322 	(g3703,g33611);
	dff 	XG1323 	(g1559,g25638);
	dff 	XG1324 	(g943,g34728);
	dff 	XG1325 	(g411,g29222);
	dff 	XG1326 	(g3953,g30449);
	dff 	XG1327 	(g3068,g25643);
	dff 	XG1328 	(g2704,g34608);
	dff 	XG1329 	(g6035,g24345);
	dff 	XG1330 	(g6082,g31922);
	dff 	XG1331 	(g49,g34994);
	dff 	XG1332 	(g1300,g25635);
	dff 	XG1333 	(g4057,g25686);
	dff 	XG1334 	(g5200,g30461);
	dff 	XG1335 	(g4843,g34466);
	dff 	XG1336 	(g5046,g31901);
	dff 	XG1337 	(g2250,g29249);
	dff 	XG1338 	(g319,g26882);
	dff 	XG1339 	(g4549,g33041);
	dff 	XG1340 	(g2453,g33011);
	dff 	XG1341 	(g5841,g25734);
	dff 	XG1342 	(g5763,g28097);
	dff 	XG1343 	(g3747,g33030);
	dff 	XG1344 	(g2912,g34618);
	dff 	XG1345 	(g2357,g33010);
	dff 	XG1346 	(g164,g31864);
	dff 	XG1347 	(g4253,g34630);
	dff 	XG1348 	(g5016,g31898);
	dff 	XG1349 	(g3119,g25653);
	dff 	XG1350 	(g1351,g25632);
	dff 	XG1351 	(g1648,g32988);
	dff 	XG1352 	(g4519,g33616);
	dff 	XG1353 	(g5115,g29280);
	dff 	XG1354 	(g3352,g33609);
	dff 	XG1355 	(g6657,g30563);
	dff 	XG1356 	(g4552,g33044);
	dff 	XG1357 	(g3893,g30437);
	dff 	XG1358 	(g3211,g30412);
	dff 	XG1359 	(g929,g21725);
	dff 	XG1360 	(g5595,g30491);
	dff 	XG1361 	(g3614,g30434);
	dff 	XG1362 	(g2894,g34612);
	dff 	XG1363 	(g3125,g29259);
	dff 	XG1364 	(g3821,g25681);
	dff 	XG1365 	(g4141,g25687);
	dff 	XG1366 	(g4570,g33617);
	dff 	XG1367 	(g5272,g30479);
	dff 	XG1368 	(g2735,g29256);
	dff 	XG1369 	(g728,g28054);
	dff 	XG1370 	(g6295,g30535);
	dff 	XG1371 	(g5417,g28094);
	dff 	XG1372 	(g2661,g30385);
	dff 	XG1373 	(g1988,g30361);
	dff 	XG1374 	(g5128,g25705);
	dff 	XG1375 	(g1548,g24260);
	dff 	XG1376 	(g3106,g29257);
	dff 	XG1377 	(g4659,g34461);
	dff 	XG1378 	(g4358,g34258);
	dff 	XG1379 	(g1792,g32993);
	dff 	XG1380 	(g2084,g33992);
	dff 	XG1381 	(g3061,g28061);
	dff 	XG1382 	(g3187,g30394);
	dff 	XG1383 	(g4311,g34449);
	dff 	XG1384 	(g2583,g34019);
	dff 	XG1385 	(g3003,g21726);
	dff 	XG1386 	(g1094,g29231);
	dff 	XG1387 	(g3841,g25682);
	dff 	XG1388 	(g4284,g21897);
	dff 	XG1389 	(g3763,g28067);
	dff 	XG1390 	(g3191,g30395);
	dff 	XG1391 	(g4239,g21892);
	dff 	XG1392 	(g3391,g31885);
	dff 	XG1393 	(g4180,g4210);
	dff 	XG1394 	(g691,g28048);
	dff 	XG1395 	(g534,g34723);
	dff 	XG1396 	(g5366,g25717);
	dff 	XG1397 	(g385,g25598);
	dff 	XG1398 	(g2004,g33987);
	dff 	XG1399 	(g2527,g30380);
	dff 	XG1400 	(g5456,g5448);
	dff 	XG1401 	(g4420,g26965);
	dff 	XG1402 	(g5148,g25706);
	dff 	XG1403 	(g4507,g30458);
	dff 	XG1404 	(g5348,g24338);
	dff 	XG1405 	(g3223,g30400);
	dff 	XG1406 	(g4931,g21904);
	dff 	XG1407 	(g2970,g34623);
	dff 	XG1408 	(g5698,g24343);
	dff 	XG1409 	(g3416,g25666);
	dff 	XG1410 	(g5260,g30473);
	dff 	XG1411 	(g1521,g24252);
	dff 	XG1412 	(g3522,g33028);
	dff 	XG1413 	(g3115,g29258);
	dff 	XG1414 	(g3251,g30407);
	dff 	XG1415 	(g1,g26958);
	dff 	XG1416 	(g4628,g34457);
	dff 	XG1417 	(g1996,g33568);
	dff 	XG1418 	(g4515,g26964);
	dff 	XG1419 	(g4300,g34735);
	dff 	XG1420 	(g1724,g30352);
	dff 	XG1421 	(g1379,g33543);
	dff 	XG1422 	(g12,g30326);
	dff 	XG1423 	(g1878,g33981);
	dff 	XG1424 	(g5619,g30500);
	dff 	XG1425 	(g71,g34786);
	dff 	XG1426 	(g59,g29277);
	not 	XG1427 	(g7266,g35);
	not 	XG1428 	(I11691,g36);
	not 	XG1429 	(I13054,g6744);
	not 	XG1430 	(I13149,g6745);
	not 	XG1431 	(I13152,g6746);
	not 	XG1432 	(I13031,g6747);
	not 	XG1433 	(I12994,g6748);
	not 	XG1434 	(I13010,g6749);
	not 	XG1435 	(I13020,g6750);
	not 	XG1436 	(I13252,g6751);
	not 	XG1437 	(I12991,g6752);
	not 	XG1438 	(I12935,g6753);
	not 	XG1439 	(g9901,g84);
	not 	XG1440 	(g10108,g120);
	not 	XG1441 	(g7231,g5);
	not 	XG1442 	(g9688,g113);
	not 	XG1443 	(g9964,g126);
	not 	XG1444 	(g9820,g99);
	not 	XG1445 	(g8286,g53);
	not 	XG1446 	(g10030,g116);
	not 	XG1447 	(g9819,g92);
	not 	XG1448 	(g8456,g56);
	not 	XG1449 	(g9581,g91);
	not 	XG1450 	(g10176,g44);
	not 	XG1451 	(g8571,g57);
	not 	XG1452 	(g9902,g100);
	not 	XG1453 	(g8356,g54);
	not 	XG1454 	(g9689,g124);
	not 	XG1455 	(g9822,g125);
	not 	XG1456 	(g9748,g114);
	not 	XG1457 	(g10073,g134);
	not 	XG1458 	(g9636,g72);
	not 	XG1459 	(g9821,g115);
	not 	XG1460 	(g10109,g135);
	not 	XG1461 	(g9534,g90);
	not 	XG1462 	(g9965,g127);
	not 	XG1463 	(g9332,g64);
	not 	XG1464 	(g9686,g73);
	not 	XG1465 	(I14827,g9686);
	not 	XG1466 	(I14679,g9332);
	not 	XG1467 	(I14970,g9965);
	not 	XG1468 	(I14742,g9534);
	not 	XG1469 	(I15073,g10109);
	not 	XG1470 	(I14902,g9821);
	not 	XG1471 	(I14797,g9636);
	not 	XG1472 	(I15030,g10073);
	not 	XG1473 	(I14866,g9748);
	not 	XG1474 	(I14905,g9822);
	not 	XG1475 	(I14839,g9689);
	not 	XG1476 	(I14241,g8356);
	not 	XG1477 	(I14935,g9902);
	not 	XG1478 	(I14301,g8571);
	not 	XG1479 	(I15162,g10176);
	not 	XG1480 	(I14773,g9581);
	not 	XG1481 	(I14271,g8456);
	not 	XG1482 	(I14893,g9819);
	not 	XG1483 	(I14999,g10030);
	not 	XG1484 	(I14222,g8286);
	not 	XG1485 	(I14896,g9820);
	not 	XG1486 	(I14967,g9964);
	not 	XG1487 	(I14836,g9688);
	not 	XG1488 	(I14079,g7231);
	not 	XG1489 	(I15070,g10108);
	not 	XG1490 	(I14932,g9901);
	not 	XG1491 	(g8989,I12935);
	not 	XG1492 	(g9153,I12991);
	not 	XG1493 	(g9637,I13252);
	not 	XG1494 	(g9213,I13020);
	not 	XG1495 	(g9186,I13010);
	not 	XG1496 	(g9154,I12994);
	not 	XG1497 	(g9245,I13031);
	not 	XG1498 	(g9478,I13152);
	not 	XG1499 	(g9477,I13149);
	not 	XG1500 	(g9280,I13054);
	not 	XG1501 	(g6869,I11691);
	not 	XG1502 	(I13847,g7266);
	not 	XG1503 	(g9716,g5057);
	not 	XG1504 	(g8579,g2771);
	not 	XG1505 	(g9590,g1882);
	nand 	XG1506 	(g9629,g6466,g6462);
	not 	XG1507 	(g9574,g6462);
	not 	XG1508 	(g7379,g2299);
	not 	XG1509 	(g8626,g4040);
	not 	XG1510 	(I12666,g4040);
	not 	XG1511 	(g10154,g2547);
	not 	XG1512 	(g9480,g559);
	not 	XG1513 	(g9049,g640);
	not 	XG1514 	(I12963,g640);
	not 	XG1515 	(g9056,g3017);
	and 	XG1516 	(g7251,g392,g452);
	nand 	XG1517 	(I13109,g5813,g5808);
	and 	XG1518 	(g8530,g2907,g2902);
	not 	XG1519 	(g9413,g1744);
	nor 	XG1520 	(g9640,g1728,g1802);
	not 	XG1521 	(g7356,g1802);
	nor 	XG1522 	(g10341,g6219,g6227);
	not 	XG1523 	(g9518,g6219);
	nand 	XG1524 	(g7850,g807,g554);
	not 	XG1525 	(I12135,g807);
	not 	XG1526 	(g8899,g807);
	not 	XG1527 	(I18700,g6027);
	nand 	XG1528 	(g9246,g812,g847);
	not 	XG1529 	(g9086,g847);
	not 	XG1530 	(g10274,g976);
	not 	XG1531 	(g6818,g976);
	or 	XG1532 	(g7673,g4172,g4153);
	not 	XG1533 	(I12861,g4372);
	not 	XG1534 	(g6958,g4372);
	not 	XG1535 	(g8021,g3512);
	not 	XG1536 	(g8770,g749);
	not 	XG1537 	(I12109,g749);
	not 	XG1538 	(g8218,g3490);
	nand 	XG1539 	(g10185,g6005,g5983,g6012,g5969);
	not 	XG1540 	(g7395,g6005);
	not 	XG1541 	(I15190,g6005);
	nand 	XG1542 	(I12840,g4235,g4222);
	or 	XG1543 	(I12902,g4226,g4229,g4232,g4235);
	not 	XG1544 	(I12899,g4232);
	not 	XG1545 	(g9250,g1600);
	not 	XG1546 	(g9970,g1714);
	not 	XG1547 	(I16606,g3649);
	not 	XG1548 	(I17852,g3625);
	not 	XG1549 	(g9916,g3625);
	not 	XG1550 	(g7964,g3155);
	nand 	XG1551 	(g9177,g3401,g3355);
	not 	XG1552 	(g9060,g3355);
	not 	XG1553 	(g10261,g4555);
	not 	XG1554 	(g8733,g3698);
	not 	XG1555 	(g9456,g6073);
	not 	XG1556 	(g9283,g1736);
	not 	XG1557 	(g10199,g1968);
	not 	XG1558 	(g7785,g4621);
	nor 	XG1559 	(g10205,g2255,g2389,g2523,g2657);
	nand 	XG1560 	(g10160,g5659,g5637,g5666,g5623);
	not 	XG1561 	(I15144,g5659);
	not 	XG1562 	(g7344,g5659);
	not 	XG1563 	(g6804,g490);
	not 	XG1564 	(g7537,g311);
	not 	XG1565 	(g7297,g6069);
	not 	XG1566 	(I12016,g772);
	not 	XG1567 	(g8859,g772);
	not 	XG1568 	(g9959,g6177);
	not 	XG1569 	(I18734,g6373);
	not 	XG1570 	(g8011,g3167);
	not 	XG1571 	(I13723,g3167);
	not 	XG1572 	(g8479,g3057);
	nand 	XG1573 	(I12372,g3462,g3457);
	not 	XG1574 	(g8068,g3457);
	nand 	XG1575 	(g8632,g1500,g1514);
	or 	XG1576 	(I12611,g1333,g1582,g1500);
	and 	XG1577 	(g10034,g1500,g1521);
	and 	XG1578 	(g9968,g1500,g1339);
	not 	XG1579 	(g7947,g1500);
	not 	XG1580 	(I12314,g1500);
	not 	XG1581 	(g8138,g1500);
	not 	XG1582 	(g7557,g1500);
	not 	XG1583 	(g7535,g1500);
	not 	XG1584 	(g9490,g2563);
	nor 	XG1585 	(g8131,g4793,g4801,g4776);
	not 	XG1586 	(g7928,g4776);
	nand 	XG1587 	(I11824,g4601,g4593);
	nand 	XG1588 	(g7227,g4593,g4584);
	not 	XG1589 	(g7163,g4593);
	not 	XG1590 	(g7072,g6199);
	not 	XG1591 	(g9339,g2295);
	nand 	XG1592 	(I12096,g1322,g1339);
	not 	XG1593 	(g7778,g1339);
	nor 	XG1594 	(g10266,g5180,g5188);
	not 	XG1595 	(g9300,g5180);
	not 	XG1596 	(g7518,g1024);
	nand 	XG1597 	(g8967,g4258,g4264);
	not 	XG1598 	(g8914,g4264);
	not 	XG1599 	(g8830,g767);
	not 	XG1600 	(I12003,g767);
	not 	XG1601 	(g7049,g5853);
	not 	XG1602 	(I16168,g3321);
	not 	XG1603 	(I18066,g3317);
	nand 	XG1604 	(I13509,g2093,g2089);
	not 	XG1605 	(g6994,g4933);
	and 	XG1606 	(g8234,g4521,g4515);
	not 	XG1607 	(g7235,g4521);
	not 	XG1608 	(g7162,g4521);
	not 	XG1609 	(g7026,g5507);
	nand 	XG1610 	(g8728,g3654,g3632,g3661,g3618);
	not 	XG1611 	(g9713,g3618);
	not 	XG1612 	(I17819,g3618);
	not 	XG1613 	(g8458,g294);
	not 	XG1614 	(I13240,g5794);
	not 	XG1615 	(g9618,g5794);
	not 	XG1616 	(g9742,g6144);
	not 	XG1617 	(I13317,g6144);
	nand 	XG1618 	(I12401,g3813,g3808);
	not 	XG1619 	(I12061,g562);
	not 	XG1620 	(g10032,g562);
	not 	XG1621 	(I12159,g608);
	not 	XG1622 	(g8945,g608);
	nor 	XG1623 	(g7661,g1205,g1221,g1216,g1211);
	and 	XG1624 	(g7918,g1087,g1205);
	not 	XG1625 	(g9174,g1205);
	not 	XG1626 	(g7851,g921);
	and 	XG1627 	(g7696,g2950,g2955);
	not 	XG1628 	(g6800,g203);
	not 	XG1629 	(g9397,g6088);
	not 	XG1630 	(g7868,g1099);
	nor 	XG1631 	(g9664,g4836,g4864,g4871,g4878);
	nand 	XG1632 	(g7846,g4878,g4843);
	not 	XG1633 	(g7991,g4878);
	not 	XG1634 	(g7840,g4878);
	not 	XG1635 	(g7521,g5630);
	not 	XG1636 	(I18555,g5630);
	not 	XG1637 	(I18509,g5623);
	not 	XG1638 	(g7470,g5623);
	nand 	XG1639 	(g9591,g1894,g1926);
	not 	XG1640 	(g8302,g1926);
	not 	XG1641 	(g9462,g6215);
	not 	XG1642 	(I12199,g6215);
	not 	XG1643 	(g8575,g291);
	nor 	XG1644 	(g9602,g4646,g4674,g4681,g4688);
	not 	XG1645 	(g7788,g4674);
	not 	XG1646 	(I15208,g637);
	not 	XG1647 	(g7496,g5969);
	not 	XG1648 	(I18560,g5969);
	not 	XG1649 	(I18728,g6012);
	not 	XG1650 	(g7471,g6012);
	nor 	XG1651 	(g9694,g1862,g1936);
	not 	XG1652 	(g7322,g1862);
	not 	XG1653 	(g8898,g676);
	not 	XG1654 	(g9220,g843);
	not 	XG1655 	(g7655,g4332);
	not 	XG1656 	(I12927,g4332);
	not 	XG1657 	(g9985,g4332);
	or 	XG1658 	(g7932,g4153,g4072);
	not 	XG1659 	(g7437,g5666);
	not 	XG1660 	(I18694,g5666);
	not 	XG1661 	(I16795,g5637);
	not 	XG1662 	(g7394,g5637);
	not 	XG1663 	(g10050,g6336);
	not 	XG1664 	(g7087,g6336);
	not 	XG1665 	(g9162,g622);
	not 	XG1666 	(I12086,g622);
	not 	XG1667 	(g7985,g3506);
	not 	XG1668 	(g7132,g4558);
	not 	XG1669 	(g7187,g6065);
	not 	XG1670 	(g7563,g6322);
	not 	XG1671 	(I18662,g6322);
	nand 	XG1672 	(g10207,g6351,g6329,g6358,g6315);
	not 	XG1673 	(g7513,g6315);
	not 	XG1674 	(I18614,g6315);
	nand 	XG1675 	(I12344,g3111,g3106);
	not 	XG1676 	(I13694,g117);
	not 	XG1677 	(I11685,g117);
	not 	XG1678 	(g10084,g2837);
	or 	XG1679 	(g7404,g939,g933);
	not 	XG1680 	(g8608,g278);
	not 	XG1681 	(g10222,g4492);
	not 	XG1682 	(I11753,g4492);
	not 	XG1683 	(g7809,g4864);
	not 	XG1684 	(g7548,g1036);
	nand 	XG1685 	(g9663,g4646,g128);
	nand 	XG1686 	(g8803,g4646,g128);
	not 	XG1687 	(g7017,g128);
	not 	XG1688 	(I13684,g128);
	and 	XG1689 	(g9967,g1157,g1178);
	not 	XG1690 	(g7715,g1178);
	not 	XG1691 	(g10074,g718);
	not 	XG1692 	(g10002,g6195);
	nand 	XG1693 	(I12203,g1135,g1094);
	not 	XG1694 	(g7069,g6137);
	not 	XG1695 	(I11801,g6395);
	not 	XG1696 	(g10169,g6395);
	not 	XG1697 	(g8155,g3380);
	not 	XG1698 	(I13360,g5343);
	not 	XG1699 	(g9856,g5343);
	not 	XG1700 	(g6808,g554);
	not 	XG1701 	(I12144,g554);
	not 	XG1702 	(g8951,g554);
	not 	XG1703 	(g6803,g496);
	not 	XG1704 	(g6926,g3853);
	not 	XG1705 	(g9671,g5134);
	not 	XG1706 	(g9011,g1422);
	not 	XG1707 	(I18337,g1422);
	not 	XG1708 	(I18297,g1418);
	not 	XG1709 	(g8955,g1418);
	not 	XG1710 	(I12523,g3794);
	not 	XG1711 	(g8345,g3794);
	nand 	XG1712 	(g9654,g2453,g2485);
	not 	XG1713 	(g8373,g2485);
	not 	XG1714 	(g7301,g925);
	not 	XG1715 	(I12415,g48);
	not 	XG1716 	(I16328,g878);
	not 	XG1717 	(I16417,g875);
	or 	XG1718 	(g8904,g1798,g1779);
	not 	XG1719 	(g7666,g4076);
	and 	XG1720 	(g8690,g2936,g2941);
	not 	XG1721 	(g8681,g763);
	not 	XG1722 	(I11992,g763);
	and 	XG1723 	(g7685,g4375,g4382);
	not 	XG1724 	(g7495,g4375);
	not 	XG1725 	(g7259,g4375);
	nand 	XG1726 	(g8889,g4871,g3684);
	nand 	XG1727 	(g9852,g4871,g3684);
	not 	XG1728 	(g7828,g4871);
	not 	XG1729 	(I12013,g590);
	not 	XG1730 	(g8851,g590);
	not 	XG1731 	(I15732,g6692);
	not 	XG1732 	(g7591,g6668);
	not 	XG1733 	(I18709,g6668);
	not 	XG1734 	(g10043,g1632);
	nand 	XG1735 	(g10124,g5313,g5290,g5320,g5276);
	not 	XG1736 	(g7296,g5313);
	not 	XG1737 	(I15102,g5313);
	not 	XG1738 	(g8438,g3100);
	not 	XG1739 	(g8216,g3092);
	not 	XG1740 	(I12451,g3092);
	not 	XG1741 	(g7876,g1495);
	not 	XG1742 	(g10058,g6497);
	not 	XG1743 	(I13374,g6490);
	not 	XG1744 	(g9818,g6490);
	nand 	XG1745 	(I12217,g1478,g1437);
	nand 	XG1746 	(I13139,g6159,g6154);
	not 	XG1747 	(g9460,g6154);
	not 	XG1748 	(g8091,g1579);
	not 	XG1749 	(I13892,g1576);
	not 	XG1750 	(g9639,g1752);
	not 	XG1751 	(g8249,g1917);
	not 	XG1752 	(I12089,g744);
	not 	XG1753 	(g8745,g744);
	not 	XG1754 	(g7975,g3040);
	not 	XG1755 	(g8673,g4737);
	not 	XG1756 	(g8133,g4809);
	not 	XG1757 	(I12411,g4809);
	not 	XG1758 	(g6900,g3440);
	nand 	XG1759 	(g8751,g4005,g3983,g4012,g3969);
	not 	XG1760 	(g9771,g3969);
	not 	XG1761 	(I17857,g3969);
	not 	XG1762 	(I17999,g4012);
	not 	XG1763 	(g9714,g4012);
	not 	XG1764 	(g7886,g1442);
	not 	XG1765 	(g10159,g4477);
	not 	XG1766 	(I13875,g1233);
	not 	XG1767 	(g7285,g4643);
	not 	XG1768 	(I16847,g6329);
	not 	XG1769 	(g7472,g6329);
	not 	XG1770 	(I15238,g6351);
	not 	XG1771 	(g7439,g6351);
	not 	XG1772 	(g8381,g2610);
	not 	XG1773 	(g7002,g5160);
	nand 	XG1774 	(g7167,g5406,g5360);
	not 	XG1775 	(g7138,g5360);
	nand 	XG1776 	(I12261,g1448,g1454);
	not 	XG1777 	(g7619,g1296);
	not 	XG1778 	(g6873,g3151);
	not 	XG1779 	(I13581,g6727);
	not 	XG1780 	(g10102,g6727);
	nor 	XG1781 	(g8906,g3522,g3530);
	not 	XG1782 	(g8165,g3530);
	not 	XG1783 	(g6990,g4742);
	not 	XG1784 	(g7670,g4104);
	nand 	XG1785 	(I13065,g4304,g4308);
	not 	XG1786 	(g9252,g4304);
	not 	XG1787 	(I13037,g4304);
	not 	XG1788 	(g9648,g2177);
	nor 	XG1789 	(g9015,g3010,g3050);
	not 	XG1790 	(g8388,g3010);
	not 	XG1791 	(I12336,g52);
	not 	XG1792 	(g6987,g4754);
	nor 	XG1793 	(g9700,g2287,g2361);
	not 	XG1794 	(g7335,g2287);
	not 	XG1795 	(g9018,g4273);
	not 	XG1796 	(I11726,g4273);
	not 	XG1797 	(g6830,g1389);
	not 	XG1798 	(g8002,g1389);
	not 	XG1799 	(g9691,g1706);
	not 	XG1800 	(g9510,g5835);
	nor 	XG1801 	(g7304,g1171,g1183);
	nand 	XG1802 	(g8609,g1157,g1171);
	not 	XG1803 	(g8407,g1171);
	not 	XG1804 	(g8964,g4269);
	not 	XG1805 	(g9832,g2399);
	not 	XG1806 	(g9360,g3372);
	nor 	XG1807 	(g8177,g4983,g4991,g4966);
	not 	XG1808 	(g9064,g4983);
	not 	XG1809 	(g9661,g3661);
	not 	XG1810 	(I17964,g3661);
	not 	XG1811 	(I12735,g4572);
	not 	XG1812 	(g8217,g3143);
	not 	XG1813 	(g6874,g3143);
	not 	XG1814 	(g8663,g3343);
	nand 	XG1815 	(I13729,g4537,g4534);
	nand 	XG1816 	(g7228,g6444,g6398);
	not 	XG1817 	(g7191,g6398);
	not 	XG1818 	(g8715,g4927);
	not 	XG1819 	(g10180,g2259);
	not 	XG1820 	(g8686,g2819);
	not 	XG1821 	(I11903,g4414);
	not 	XG1822 	(g7258,g4414);
	not 	XG1823 	(g9887,g5802);
	not 	XG1824 	(g9333,g417);
	not 	XG1825 	(g9903,g681);
	not 	XG1826 	(I12997,g351);
	or 	XG1827 	(g7834,g2946,g2886);
	not 	XG1828 	(g8281,g3494);
	not 	XG1829 	(g6904,g3494);
	not 	XG1830 	(g9239,g5511);
	not 	XG1831 	(g8070,g3518);
	not 	XG1832 	(I13744,g3518);
	not 	XG1833 	(g7267,g1604);
	nand 	XG1834 	(g9724,g5084,g5092);
	not 	XG1835 	(g9669,g5092);
	nand 	XG1836 	(g8847,g4681,g4831);
	nand 	XG1837 	(g9775,g4681,g4831);
	not 	XG1838 	(g7063,g4831);
	and 	XG1839 	(g7469,g4438,g4382);
	not 	XG1840 	(g7289,g4382);
	not 	XG1841 	(g10191,g6386);
	not 	XG1842 	(g7410,g2008);
	not 	XG1843 	(g8836,g736);
	not 	XG1844 	(g9905,g802);
	not 	XG1845 	(I14563,g802);
	or 	XG1846 	(g8679,g199,g222);
	nand 	XG1847 	(g9092,g3050,g3004);
	not 	XG1848 	(g8340,g3050);
	not 	XG1849 	(g9733,g5736);
	not 	XG1850 	(g7913,g1052);
	not 	XG1851 	(I12538,g58);
	not 	XG1852 	(g10152,g2122);
	not 	XG1853 	(g7424,g2465);
	not 	XG1854 	(g7092,g6483);
	nor 	XG1855 	(g8720,g365,g358);
	and 	XG1856 	(g8721,g365,g376,g385);
	not 	XG1857 	(I12719,g365);
	nand 	XG1858 	(g7836,g4688,g4653);
	nand 	XG1859 	(g7690,g4653,g4659,g4669);
	not 	XG1860 	(g8606,g4653);
	nor 	XG1861 	(g8864,g3171,g3179);
	not 	XG1862 	(g8107,g3179);
	not 	XG1863 	(g7275,g1728);
	not 	XG1864 	(g7423,g2433);
	not 	XG1865 	(g8228,g3835);
	not 	XG1866 	(g9620,g6187);
	not 	XG1867 	(g6820,g1070);
	not 	XG1868 	(g7750,g1070);
	and 	XG1869 	(g7777,g817,g822,g723);
	not 	XG1870 	(g7216,g822);
	not 	XG1871 	(I16770,g6023);
	not 	XG1872 	(g7443,g914);
	not 	XG1873 	(I18600,g5335);
	not 	XG1874 	(I11701,g4164);
	or 	XG1875 	(g9483,g969,g1008);
	not 	XG1876 	(g7903,g969);
	not 	XG1877 	(g8639,g2807);
	nand 	XG1878 	(g9442,g5428,g5424);
	not 	XG1879 	(g9379,g5424);
	not 	XG1880 	(g8700,g4054);
	not 	XG1881 	(I11716,g4054);
	not 	XG1882 	(g9684,g6191);
	not 	XG1883 	(g7073,g6191);
	not 	XG1884 	(g9989,g5077);
	not 	XG1885 	(I12176,g5523);
	not 	XG1886 	(g9311,g5523);
	not 	XG1887 	(I17938,g3676);
	nor 	XG1888 	(g8086,g182,g174,g168);
	not 	XG1889 	(g9969,g1682);
	nor 	XG1890 	(g7499,g355,g333);
	not 	XG1891 	(g9050,g1087);
	not 	XG1892 	(g8654,g1087);
	not 	XG1893 	(g9007,g1083);
	not 	XG1894 	(I18333,g1083);
	nand 	XG1895 	(I12240,g1105,g1111);
	not 	XG1896 	(g8267,g2342);
	not 	XG1897 	(g8565,g3802);
	not 	XG1898 	(g8659,g2815);
	not 	XG1899 	(g7400,g911);
	not 	XG1900 	(I11860,g43);
	not 	XG1901 	(I16246,g3983);
	not 	XG1902 	(g9662,g3983);
	not 	XG1903 	(g9537,g1748);
	not 	XG1904 	(g9316,g5742);
	not 	XG1905 	(g9557,g5499);
	not 	XG1906 	(g7027,g5499);
	and 	XG1907 	(g7763,g2960,g2965);
	not 	XG1908 	(g6991,g4888);
	not 	XG1909 	(g7497,g6358);
	not 	XG1910 	(I18752,g6358);
	nand 	XG1911 	(g7582,g1373,g1361);
	not 	XG1912 	(g8033,g157);
	not 	XG1913 	(g8635,g2783);
	nand 	XG1914 	(I12848,g4277,g4281);
	not 	XG1915 	(g8840,g4277);
	not 	XG1916 	(I12819,g4277);
	not 	XG1917 	(g9973,g2112);
	or 	XG1918 	(g7450,g1283,g1277);
	nor 	XG1919 	(g10123,g4297,g4294);
	not 	XG1920 	(I13623,g4294);
	not 	XG1921 	(g7438,g5983);
	not 	XG1922 	(I16821,g5983);
	not 	XG1923 	(I15837,g1459);
	not 	XG1924 	(g8301,g1399);
	not 	XG1925 	(I19837,g1399);
	not 	XG1926 	(I12123,g758);
	not 	XG1927 	(g8651,g758);
	nor 	XG1928 	(g7158,g5712,g5752);
	not 	XG1929 	(g9807,g5712);
	not 	XG1930 	(g6954,g4138);
	not 	XG1931 	(g7202,g4639);
	not 	XG1932 	(g7096,g6537);
	not 	XG1933 	(g9745,g6537);
	not 	XG1934 	(I12608,g1582);
	not 	XG1935 	(g8443,g3736);
	and 	XG1936 	(g9217,g626,g632);
	not 	XG1937 	(g6814,g632);
	not 	XG1938 	(I12120,g632);
	not 	XG1939 	(g9000,g632);
	not 	XG1940 	(I12577,g1227);
	not 	XG1941 	(I15536,g1227);
	not 	XG1942 	(g8442,g3476);
	or 	XG1943 	(g8863,g1664,g1644);
	not 	XG1944 	(I11655,g1246);
	not 	XG1945 	(g8056,g1246);
	nand 	XG1946 	(g9954,g6120,g6128);
	not 	XG1947 	(g9889,g6128);
	nand 	XG1948 	(I13382,g246,g269);
	not 	XG1949 	(g8296,g246);
	not 	XG1950 	(g8756,g4049);
	not 	XG1951 	(g7261,g4449);
	not 	XG1952 	(I11908,g4449);
	or 	XG1953 	(g7764,g2932,g2999);
	not 	XG1954 	(g6957,g2932);
	not 	XG1955 	(I12749,g4575);
	not 	XG1956 	(g6989,g4575);
	not 	XG1957 	(g7636,g4098);
	not 	XG1958 	(I12805,g4098);
	not 	XG1959 	(I12360,g528);
	not 	XG1960 	(g8046,g528);
	nand 	XG1961 	(g9800,g5428,g5436);
	not 	XG1962 	(g9730,g5436);
	not 	XG1963 	(I11632,g16);
	not 	XG1964 	(g10106,g16);
	not 	XG1965 	(g8154,g3139);
	not 	XG1966 	(I13637,g102);
	nand 	XG1967 	(I13749,g4584,g4608);
	not 	XG1968 	(g10275,g4584);
	not 	XG1969 	(g8297,g142);
	not 	XG1970 	(I16713,g5331);
	not 	XG1971 	(g9888,g5831);
	nand 	XG1972 	(I13442,g239,g262);
	not 	XG1973 	(g8363,g239);
	not 	XG1974 	(g9223,g1216);
	not 	XG1975 	(g9932,g5805);
	not 	XG1976 	(g9681,g5798);
	not 	XG1977 	(I13276,g5798);
	nor 	XG1978 	(g10338,g5022,g5062);
	not 	XG1979 	(g9670,g5022);
	not 	XG1980 	(I18107,g4019);
	not 	XG1981 	(I16639,g4000);
	nand 	XG1982 	(g7549,g1030,g1018);
	not 	XG1983 	(I16181,g3672);
	not 	XG1984 	(I18092,g3668);
	and 	XG1985 	(g7948,g1430,g1548);
	not 	XG1986 	(g8685,g1430);
	not 	XG1987 	(g9091,g1430);
	not 	XG1988 	(g9051,g1426);
	not 	XG1989 	(I18360,g1426);
	not 	XG1990 	(g7293,g4452);
	not 	XG1991 	(I11896,g4446);
	not 	XG1992 	(g7246,g4446);
	not 	XG1993 	(g10038,g2241);
	nor 	XG1994 	(g7675,g1548,g1564,g1559,g1554);
	not 	XG1995 	(g9226,g1564);
	not 	XG1996 	(g9958,g6148);
	not 	XG1997 	(I13280,g6140);
	not 	XG1998 	(g9683,g6140);
	not 	XG1999 	(I13287,g110);
	not 	XG2000 	(I16357,g884);
	not 	XG2001 	(I16345,g881);
	not 	XG2002 	(g8075,g3742);
	not 	XG2003 	(g8457,g225);
	not 	XG2004 	(g10184,g4486);
	nor 	XG2005 	(g10312,g5873,g5881);
	not 	XG2006 	(g9451,g5873);
	not 	XG2007 	(g9253,g5037);
	nand 	XG2008 	(g9595,g2319,g2351);
	not 	XG2009 	(g8211,g2319);
	not 	XG2010 	(g9500,g5495);
	not 	XG2011 	(I14619,g4185);
	not 	XG2012 	(g6846,g2152);
	not 	XG2013 	(g9392,g5869);
	not 	XG2014 	(I12189,g5869);
	not 	XG2015 	(g7170,g5719);
	not 	XG2016 	(I11665,g1589);
	not 	XG2017 	(g8092,g1589);
	nand 	XG2018 	(g7184,g5752,g5706);
	not 	XG2019 	(g9739,g5752);
	and 	XG2020 	(g7804,g2970,g2975);
	not 	XG2021 	(g9816,g6167);
	not 	XG2022 	(I14424,g4005);
	not 	XG2023 	(g9601,g4005);
	not 	XG2024 	(g7462,g2599);
	nor 	XG2025 	(g9100,g3712,g3752);
	not 	XG2026 	(g8507,g3712);
	not 	XG2027 	(g9206,g5164);
	nor 	XG2028 	(g7601,g1333,g1322);
	not 	XG2029 	(g8240,g1333);
	not 	XG2030 	(g7995,g153);
	not 	XG2031 	(g9407,g6549);
	not 	XG2032 	(I12746,g4087);
	not 	XG2033 	(g7697,g4087);
	not 	XG2034 	(g7892,g4801);
	nand 	XG2035 	(g9509,g5774,g5770);
	not 	XG2036 	(g9449,g5770);
	not 	XG2037 	(g7517,g962);
	not 	XG2038 	(I11835,g101);
	not 	XG2039 	(I12893,g4226);
	or 	XG2040 	(I12903,g4213,g4216,g4219,g4222);
	not 	XG2041 	(I12837,g4222);
	not 	XG2042 	(I12572,g51);
	not 	XG2043 	(g8734,g4045);
	nand 	XG2044 	(I12277,g1472,g1467);
	not 	XG2045 	(g10158,g2461);
	not 	XG2046 	(g7157,g5706);
	not 	XG2047 	(I11682,g2756);
	not 	XG2048 	(g9978,g2756);
	not 	XG2049 	(g9992,g5990);
	not 	XG2050 	(g7064,g5990);
	not 	XG2051 	(g7446,g1256);
	not 	XG2052 	(g7134,g5029);
	not 	XG2053 	(g9962,g6519);
	not 	XG2054 	(g7824,g4169);
	not 	XG2055 	(g10036,g1816);
	not 	XG2056 	(g8497,g3436);
	not 	XG2057 	(g9880,g5787);
	not 	XG2058 	(g6997,g4578);
	not 	XG2059 	(I12793,g4578);
	not 	XG2060 	(g10308,g4459);
	not 	XG2061 	(g8566,g3831);
	nand 	XG2062 	(I13518,g2518,g2514);
	not 	XG2063 	(g8531,g3288);
	not 	XG2064 	(g6895,g3288);
	not 	XG2065 	(g9913,g2403);
	and 	XG2066 	(g7511,g2130,g2138,g2145);
	not 	XG2067 	(g6841,g2145);
	not 	XG2068 	(g10150,g1700);
	not 	XG2069 	(g9158,g513);
	not 	XG2070 	(g10119,g2841);
	not 	XG2071 	(g9853,g5297);
	not 	XG2072 	(g7018,g5297);
	not 	XG2073 	(g8592,g3805);
	not 	XG2074 	(I12563,g3798);
	not 	XG2075 	(g8399,g3798);
	not 	XG2076 	(g9657,g2763);
	not 	XG2077 	(g9030,g4793);
	not 	XG2078 	(g7597,g952);
	not 	XG2079 	(g7577,g1263);
	not 	XG2080 	(g10079,g1950);
	not 	XG2081 	(g9729,g5138);
	not 	XG2082 	(g9594,g2307);
	not 	XG2083 	(g9728,g5109);
	not 	XG2084 	(I13166,g5101);
	not 	XG2085 	(g9498,g5101);
	not 	XG2086 	(g7046,g5791);
	not 	XG2087 	(g8650,g4664);
	or 	XG2088 	(g8905,g2223,g2204);
	not 	XG2089 	(g9390,g5808);
	not 	XG2090 	(g9644,g2016);
	not 	XG2091 	(g9933,g5759);
	nor 	XG2092 	(g8958,g3873,g3881);
	not 	XG2093 	(g8172,g3873);
	not 	XG2094 	(g9600,g3632);
	not 	XG2095 	(I16217,g3632);
	not 	XG2096 	(g9552,g3654);
	not 	XG2097 	(I14395,g3654);
	not 	XG2098 	(g9760,g2315);
	or 	XG2099 	(g9012,g2066,g2047);
	not 	XG2100 	(g8125,g3869);
	not 	XG2101 	(I11820,g3869);
	not 	XG2102 	(g9180,g3719);
	not 	XG2103 	(I12355,g46);
	nand 	XG2104 	(g9203,g3752,g3706);
	not 	XG2105 	(g8449,g3752);
	or 	XG2106 	(I12782,g4200,g4197,g4194,g4188);
	not 	XG2107 	(I12761,g4188);
	not 	XG2108 	(I14450,g4191);
	not 	XG2109 	(I12654,g1585);
	not 	XG2110 	(g8364,g1585);
	not 	XG2111 	(I12605,g1570);
	not 	XG2112 	(I15542,g1570);
	nand 	XG2113 	(I11877,g4430,g4388);
	not 	XG2114 	(I12887,g4216);
	not 	XG2115 	(I12884,g4213);
	not 	XG2116 	(g10183,g2595);
	not 	XG2117 	(g9976,g2537);
	not 	XG2118 	(I13708,g136);
	not 	XG2119 	(g10139,g136);
	not 	XG2120 	(g7149,g4564);
	not 	XG2121 	(I11743,g4564);
	not 	XG2122 	(g8539,g3454);
	not 	XG2123 	(g8343,g3447);
	not 	XG2124 	(I12519,g3447);
	not 	XG2125 	(g8764,g4826);
	not 	XG2126 	(g8713,g4826);
	not 	XG2127 	(g7086,g4826);
	nand 	XG2128 	(g8227,g3774,g3770);
	not 	XG2129 	(g8170,g3770);
	nand 	XG2130 	(I13497,g232,g255);
	not 	XG2131 	(g8406,g232);
	not 	XG2132 	(g7095,g6545);
	not 	XG2133 	(g10153,g2417);
	not 	XG2134 	(g6848,g2417);
	not 	XG2135 	(g7315,g1772);
	not 	XG2136 	(g9229,g5052);
	not 	XG2137 	(g9616,g5452);
	not 	XG2138 	(I13236,g5452);
	not 	XG2139 	(g9753,g1890);
	nor 	XG2140 	(g9835,g2555,g2629);
	not 	XG2141 	(g7490,g2629);
	not 	XG2142 	(I12103,g572);
	not 	XG2143 	(g8766,g572);
	not 	XG2144 	(g7680,g4108);
	nor 	XG2145 	(g7567,g990,g979);
	or 	XG2146 	(I12583,g990,g1239,g1157);
	not 	XG2147 	(g8186,g990);
	not 	XG2148 	(I12580,g1239);
	not 	XG2149 	(g10197,g31);
	not 	XG2150 	(I11626,g31);
	not 	XG2151 	(g8538,g3412);
	not 	XG2152 	(I12333,g45);
	not 	XG2153 	(I15036,g799);
	not 	XG2154 	(g9099,g3706);
	not 	XG2155 	(g8623,g3990);
	not 	XG2156 	(g6941,g3990);
	not 	XG2157 	(g9434,g5385);
	not 	XG2158 	(g9511,g5881);
	not 	XG2159 	(g6840,g1992);
	not 	XG2160 	(g10151,g1992);
	not 	XG2161 	(g8097,g3029);
	not 	XG2162 	(g8059,g3171);
	not 	XG2163 	(g8558,g3787);
	not 	XG2164 	(g7197,g812);
	nand 	XG2165 	(g9334,g832,g827);
	not 	XG2166 	(g7118,g832);
	not 	XG2167 	(g7765,g4165);
	nand 	XG2168 	(g8691,g3303,g3281,g3310,g3267);
	not 	XG2169 	(g9551,g3281);
	not 	XG2170 	(I16193,g3281);
	not 	XG2171 	(I14365,g3303);
	not 	XG2172 	(g9496,g3303);
	not 	XG2173 	(g6917,g3684);
	not 	XG2174 	(g6918,g3639);
	not 	XG2175 	(g8584,g3639);
	not 	XG2176 	(I18795,g5327);
	not 	XG2177 	(I12618,g3338);
	not 	XG2178 	(g8534,g3338);
	nor 	XG2179 	(g7139,g5366,g5406);
	not 	XG2180 	(g9678,g5406);
	not 	XG2181 	(g6923,g3791);
	not 	XG2182 	(g8136,g269);
	not 	XG2183 	(g10166,g6040);
	and 	XG2184 	(g7396,g441,g392);
	not 	XG2185 	(I13202,g5105);
	not 	XG2186 	(g9554,g5105);
	not 	XG2187 	(g8123,g3808);
	not 	XG2188 	(g10072,g9);
	not 	XG2189 	(I11635,g9);
	not 	XG2190 	(g8593,g3759);
	not 	XG2191 	(I11737,g4467);
	not 	XG2192 	(I12758,g4093);
	not 	XG2193 	(g7733,g4093);
	nand 	XG2194 	(g9538,g1760,g1792);
	not 	XG2195 	(g8146,g1760);
	not 	XG2196 	(g10000,g6151);
	not 	XG2197 	(g8287,g160);
	not 	XG2198 	(g7023,g5445);
	not 	XG2199 	(g7153,g5373);
	not 	XG2200 	(g10081,g2279);
	not 	XG2201 	(g8541,g3498);
	not 	XG2202 	(I12117,g586);
	not 	XG2203 	(g10262,g586);
	not 	XG2204 	(I16401,g869);
	not 	XG2205 	(I16391,g859);
	nand 	XG2206 	(g9705,g2587,g2619);
	not 	XG2207 	(g8418,g2619);
	not 	XG2208 	(g8462,g1183);
	not 	XG2209 	(g9337,g1608);
	not 	XG2210 	(I12767,g4197);
	not 	XG2211 	(I12764,g4194);
	not 	XG2212 	(g7512,g5283);
	not 	XG2213 	(I18504,g5283);
	not 	XG2214 	(g7436,g5276);
	not 	XG2215 	(I18460,g5276);
	nand 	XG2216 	(I13564,g2652,g2648);
	not 	XG2217 	(g10040,g2652);
	not 	XG2218 	(g9861,g5459);
	not 	XG2219 	(g10086,g2193);
	not 	XG2220 	(g10203,g2393);
	not 	XG2221 	(g10096,g5767);
	not 	XG2222 	(g10110,g661);
	nor 	XG2223 	(g10281,g5527,g5535);
	not 	XG2224 	(g9444,g5535);
	not 	XG2225 	(g9152,g2834);
	nand 	XG2226 	(g8163,g3423,g3419);
	not 	XG2227 	(g8112,g3419);
	not 	XG2228 	(g7845,g1146);
	or 	XG2229 	(g9055,g2625,g2606);
	not 	XG2230 	(g9073,g150);
	nor 	XG2231 	(g10179,g1696,g1830,g1964,g2098);
	not 	XG2232 	(g9472,g6555);
	not 	XG2233 	(g8390,g3385);
	not 	XG2234 	(g8229,g3881);
	not 	XG2235 	(g8397,g3470);
	not 	XG2236 	(g9187,g518);
	not 	XG2237 	(g8005,g3025);
	or 	XG2238 	(g9535,g538,g209);
	not 	XG2239 	(g10136,g6113);
	not 	XG2240 	(g9374,g5188);
	not 	XG2241 	(I13424,g5689);
	not 	XG2242 	(g9927,g5689);
	not 	XG2243 	(I15824,g1116);
	not 	XG2244 	(I19818,g1056);
	not 	XG2245 	(g8239,g1056);
	nor 	XG2246 	(g8182,g392,g405);
	nand 	XG2247 	(I12468,g392,g405);
	not 	XG2248 	(g8037,g405);
	not 	XG2249 	(g10026,g6494);
	not 	XG2250 	(g9744,g6486);
	not 	XG2251 	(I13321,g6486);
	not 	XG2252 	(g8672,g4669);
	not 	XG2253 	(g6985,g4669);
	not 	XG2254 	(g9439,g5428);
	not 	XG2255 	(g9070,g5428);
	nand 	XG2256 	(I12074,g979,g996);
	and 	XG2257 	(g9906,g1157,g996);
	not 	XG2258 	(g7749,g996);
	not 	XG2259 	(g6982,g4531);
	not 	XG2260 	(g6986,g4743);
	nand 	XG2261 	(g8292,g215,g218);
	not 	XG2262 	(I12503,g215);
	not 	XG2263 	(g7232,g4411);
	not 	XG2264 	(g6831,g1413);
	not 	XG2265 	(g7779,g1413);
	not 	XG2266 	(I11750,g4474);
	not 	XG2267 	(I15663,g5308);
	not 	XG2268 	(g8426,g3045);
	not 	XG2269 	(g9900,g6);
	not 	XG2270 	(g7405,g1936);
	not 	XG2271 	(I12418,g55);
	not 	XG2272 	(g9077,g504);
	not 	XG2273 	(g8330,g2587);
	not 	XG2274 	(g9699,g2311);
	not 	XG2275 	(g6802,g468);
	not 	XG2276 	(g9556,g5448);
	not 	XG2277 	(I13206,g5448);
	not 	XG2278 	(g8669,g3767);
	not 	XG2279 	(g9808,g5827);
	not 	XG2280 	(g7970,g4688);
	not 	XG2281 	(g7827,g4688);
	nand 	XG2282 	(g9883,g5774,g5782);
	not 	XG2283 	(g9103,g5774);
	not 	XG2284 	(g9506,g5774);
	nand 	XG2285 	(I13462,g2384,g2380);
	not 	XG2286 	(g9264,g5396);
	not 	XG2287 	(g9754,g2020);
	not 	XG2288 	(I17901,g3976);
	not 	XG2289 	(g9982,g3976);
	not 	XG2290 	(I18293,g1079);
	not 	XG2291 	(g8954,g1079);
	not 	XG2292 	(g8903,g1075);
	not 	XG2293 	(I18276,g1075);
	not 	XG2294 	(g10060,g6541);
	nor 	XG2295 	(g9586,g1592,g1668);
	not 	XG2296 	(g7308,g1668);
	not 	XG2297 	(g8180,g262);
	not 	XG2298 	(g9752,g1840);
	not 	XG2299 	(I11688,g70);
	nand 	XG2300 	(I13077,g5467,g5462);
	not 	XG2301 	(g9402,g6209);
	not 	XG2302 	(I13606,g74);
	not 	XG2303 	(g7631,g74);
	not 	XG2304 	(g7343,g5290);
	not 	XG2305 	(I16762,g5290);
	not 	XG2306 	(g10033,g655);
	not 	XG2307 	(g6903,g3502);
	not 	XG2308 	(g7236,g4608);
	not 	XG2309 	(g7183,g4608);
	not 	XG2310 	(g8833,g794);
	not 	XG2311 	(I12112,g794);
	not 	XG2312 	(I16201,g4023);
	not 	XG2313 	(I13726,g4537);
	not 	XG2314 	(I12644,g3689);
	not 	XG2315 	(g8587,g3689);
	not 	XG2316 	(g9305,g5381);
	not 	XG2317 	(I18653,g5681);
	not 	XG2318 	(g9582,g703);
	not 	XG2319 	(g10047,g5421);
	not 	XG2320 	(g7441,g862);
	not 	XG2321 	(g7411,g2040);
	not 	XG2322 	(I12437,g4999);
	not 	XG2323 	(g8179,g4999);
	not 	XG2324 	(I13352,g4146);
	not 	XG2325 	(g7963,g4146);
	not 	XG2326 	(g10311,g4633);
	not 	XG2327 	(g7532,g1157);
	not 	XG2328 	(g7917,g1157);
	not 	XG2329 	(I12300,g1157);
	not 	XG2330 	(g7519,g1157);
	not 	XG2331 	(g8087,g1157);
	not 	XG2332 	(g7262,g5723);
	not 	XG2333 	(g9450,g5817);
	not 	XG2334 	(g8316,g2351);
	not 	XG2335 	(g10229,g6736);
	not 	XG2336 	(g6995,g4944);
	or 	XG2337 	(g7684,g4176,g4072);
	not 	XG2338 	(g7541,g344);
	not 	XG2339 	(I12026,g344);
	not 	XG2340 	(g7340,g4443);
	not 	XG2341 	(g8113,g3466);
	not 	XG2342 	(g9364,g5041);
	not 	XG2343 	(g9797,g5441);
	nand 	XG2344 	(I11864,g4401,g4434);
	not 	XG2345 	(g8508,g3827);
	nand 	XG2346 	(I13182,g6505,g6500);
	not 	XG2347 	(g9527,g6500);
	not 	XG2348 	(I18813,g5673);
	not 	XG2349 	(I15677,g5654);
	not 	XG2350 	(g8106,g3133);
	not 	XG2351 	(g8718,g3333);
	not 	XG2352 	(g8765,g3333);
	not 	XG2353 	(g6887,g3333);
	not 	XG2354 	(g6825,g979);
	not 	XG2355 	(g7806,g4681);
	not 	XG2356 	(g8522,g298);
	nand 	XG2357 	(g8561,g3774,g3782);
	not 	XG2358 	(g7952,g3774);
	not 	XG2359 	(g8224,g3774);
	not 	XG2360 	(g9977,g2667);
	not 	XG2361 	(g8492,g3396);
	or 	XG2362 	(I12783,g4180,g4210,g4207,g4204);
	not 	XG2363 	(I12779,g4210);
	not 	XG2364 	(I12776,g4207);
	not 	XG2365 	(g8201,g1894);
	or 	XG2366 	(g8461,g534,g301);
	not 	XG2367 	(g6809,g341);
	not 	XG2368 	(g9194,g827);
	not 	XG2369 	(g9559,g6077);
	not 	XG2370 	(g7431,g2555);
	nand 	XG2371 	(g9715,g4836,g5011);
	nand 	XG2372 	(g8829,g4836,g5011);
	not 	XG2373 	(g7109,g5011);
	not 	XG2374 	(g6799,g199);
	not 	XG2375 	(g10027,g6523);
	nor 	XG2376 	(g7352,g1514,g1526);
	not 	XG2377 	(g8526,g1526);
	not 	XG2378 	(g7224,g4601);
	nand 	XG2379 	(I12287,g1300,g1484);
	nand 	XG2380 	(g9372,g5084,g5080);
	not 	XG2381 	(g9298,g5080);
	not 	XG2382 	(g9321,g5863);
	not 	XG2383 	(I13699,g4581);
	not 	XG2384 	(g9291,g3021);
	not 	XG2385 	(g9974,g2518);
	not 	XG2386 	(g7461,g2567);
	not 	XG2387 	(g10143,g568);
	not 	XG2388 	(I12083,g568);
	not 	XG2389 	(g10190,g6044);
	nor 	XG2390 	(g7192,g6404,g6444);
	not 	XG2391 	(g9898,g6444);
	not 	XG2392 	(g9274,g5857);
	not 	XG2393 	(g9585,g1616);
	nand 	XG2394 	(g7442,g890,g896);
	not 	XG2395 	(I13718,g890);
	not 	XG2396 	(g7397,g890);
	not 	XG2397 	(g7536,g5976);
	not 	XG2398 	(I18609,g5976);
	not 	XG2399 	(g7960,g1404);
	not 	XG2400 	(g9429,g3723);
	not 	XG2401 	(g8171,g3817);
	not 	XG2402 	(I11816,g93);
	not 	XG2403 	(g8519,g287);
	not 	XG2404 	(I13094,g2724);
	not 	XG2405 	(g9839,g2724);
	nor 	XG2406 	(g10318,g22,g25);
	not 	XG2407 	(g7116,g22);
	not 	XG2408 	(g7780,g2878);
	not 	XG2409 	(g9214,g617);
	not 	XG2410 	(I12064,g617);
	not 	XG2411 	(g6827,g1277);
	not 	XG2412 	(g9899,g6513);
	not 	XG2413 	(g7564,g336);
	not 	XG2414 	(g6816,g933);
	not 	XG2415 	(g7362,g1906);
	and 	XG2416 	(g9479,g324,g305);
	not 	XG2417 	(g7523,g305);
	not 	XG2418 	(g10028,g8);
	not 	XG2419 	(g9095,g3368);
	not 	XG2420 	(I16371,g887);
	not 	XG2421 	(g7908,g4157);
	not 	XG2422 	(I13473,g4157);
	not 	XG2423 	(g6953,g4157);
	not 	XG2424 	(g10118,g2541);
	nor 	XG2425 	(g9649,g2153,g2227);
	not 	XG2426 	(g7280,g2153);
	not 	XG2427 	(g8743,g550);
	not 	XG2428 	(g8237,g255);
	nand 	XG2429 	(g8434,g3072,g3080);
	not 	XG2430 	(g8387,g3080);
	not 	XG2431 	(g8080,g3863);
	nand 	XG2432 	(I13452,g1959,g1955);
	not 	XG2433 	(g9907,g1959);
	not 	XG2434 	(g8505,g3480);
	not 	XG2435 	(I18758,g6719);
	not 	XG2436 	(I16829,g6715);
	not 	XG2437 	(I16741,g5677);
	not 	XG2438 	(g8026,g3857);
	not 	XG2439 	(g9040,g499);
	not 	XG2440 	(g9862,g5413);
	not 	XG2441 	(g7635,g1002);
	not 	XG2442 	(g8748,g776);
	not 	XG2443 	(I12033,g776);
	not 	XG2444 	(g10175,g28);
	not 	XG2445 	(I11623,g28);
	not 	XG2446 	(g8055,g1236);
	not 	XG2447 	(g8350,g4646);
	not 	XG2448 	(g8324,g2476);
	nand 	XG2449 	(g9485,g1624,g1657);
	not 	XG2450 	(g8187,g1657);
	not 	XG2451 	(g10082,g2375);
	not 	XG2452 	(I13705,g63);
	nand 	XG2453 	(g8678,g358,g376);
	nand 	XG2454 	(g8806,g385,g376,g370,g358);
	not 	XG2455 	(g8848,g358);
	not 	XG2456 	(g7475,g896);
	nand 	XG2457 	(g8500,g3423,g3431);
	not 	XG2458 	(g7926,g3423);
	not 	XG2459 	(g8160,g3423);
	not 	XG2460 	(g8631,g283);
	not 	XG2461 	(g7980,g3161);
	not 	XG2462 	(g9911,g2384);
	nor 	XG2463 	(g9061,g3361,g3401);
	not 	XG2464 	(g8441,g3361);
	nand 	XG2465 	(g10224,g6697,g6675,g6704,g6661);
	not 	XG2466 	(I16875,g6675);
	not 	XG2467 	(g7498,g6675);
	not 	XG2468 	(I15284,g6697);
	not 	XG2469 	(g7473,g6697);
	not 	XG2470 	(g6978,g4616);
	not 	XG2471 	(g10223,g4561);
	not 	XG2472 	(g9828,g2024);
	not 	XG2473 	(g8504,g3451);
	not 	XG2474 	(I12487,g3443);
	not 	XG2475 	(g8280,g3443);
	not 	XG2476 	(g8854,g613);
	not 	XG2477 	(I12046,g613);
	not 	XG2478 	(g10232,g4527);
	not 	XG2479 	(g9826,g1844);
	not 	XG2480 	(g8478,g3103);
	not 	XG2481 	(g8278,g3096);
	not 	XG2482 	(I12483,g3096);
	not 	XG2483 	(g10155,g2643);
	not 	XG2484 	(g9999,g6109);
	not 	XG2485 	(g7867,g1489);
	not 	XG2486 	(g9672,g5390);
	nand 	XG2487 	(I12544,g194,g191);
	not 	XG2488 	(g8362,g194);
	not 	XG2489 	(I12541,g194);
	not 	XG2490 	(g10181,g2551);
	not 	XG2491 	(g6849,g2551);
	not 	XG2492 	(g9779,g5156);
	nand 	XG2493 	(g8105,g3072,g3068);
	not 	XG2494 	(g8102,g3072);
	not 	XG2495 	(g7907,g3072);
	not 	XG2496 	(g8300,g1242);
	not 	XG2497 	(I12631,g1242);
	not 	XG2498 	(I12382,g47);
	not 	XG2499 	(g10133,g6049);
	not 	XG2500 	(I11793,g6049);
	not 	XG2501 	(g8334,g3034);
	not 	XG2502 	(g10039,g2273);
	not 	XG2503 	(I18845,g6711);
	nor 	XG2504 	(g7175,g6058,g6098);
	nand 	XG2505 	(g7209,g6098,g6052);
	not 	XG2506 	(g9815,g6098);
	not 	XG2507 	(g8480,g3147);
	not 	XG2508 	(g8696,g3347);
	not 	XG2509 	(g9831,g2269);
	not 	XG2510 	(I12106,g626);
	not 	XG2511 	(g9083,g626);
	not 	XG2512 	(g9491,g2729);
	not 	XG2513 	(I13124,g2729);
	not 	XG2514 	(I11777,g5357);
	not 	XG2515 	(g10044,g5357);
	not 	XG2516 	(g7898,g4991);
	not 	XG2517 	(I18825,g6019);
	not 	XG2518 	(I15697,g6000);
	nor 	XG2519 	(g8933,g4785,g4709);
	not 	XG2520 	(g8883,g4709);
	not 	XG2521 	(g6984,g4709);
	not 	XG2522 	(g9523,g6419);
	not 	XG2523 	(g7174,g6052);
	and 	XG2524 	(g8643,g2922,g2927);
	nand 	XG2525 	(g8347,g4340,g4349,g4358);
	not 	XG2526 	(I12790,g4340);
	not 	XG2527 	(I12910,g4340);
	not 	XG2528 	(I12858,g4340);
	not 	XG2529 	(I12811,g4340);
	not 	XG2530 	(g8928,g4340);
	not 	XG2531 	(I16575,g3298);
	not 	XG2532 	(g6940,g4035);
	not 	XG2533 	(g8742,g4035);
	not 	XG2534 	(g8804,g4035);
	not 	XG2535 	(g7544,g918);
	not 	XG2536 	(g8567,g4082);
	not 	XG2537 	(g10157,g2036);
	not 	XG2538 	(g8997,g577);
	not 	XG2539 	(I12132,g577);
	not 	XG2540 	(g9638,g1620);
	not 	XG2541 	(g9071,g2831);
	not 	XG2542 	(g7528,g930);
	not 	XG2543 	(g9806,g5782);
	not 	XG2544 	(g10320,g817);
	not 	XG2545 	(g7863,g1249);
	not 	XG2546 	(g9166,g837);
	not 	XG2547 	(I12141,g599);
	not 	XG2548 	(g8895,g599);
	not 	XG2549 	(g9679,g5475);
	not 	XG2550 	(I12067,g739);
	not 	XG2551 	(g8725,g739);
	not 	XG2552 	(g7110,g6682);
	not 	XG2553 	(g10099,g6682);
	not 	XG2554 	(g10001,g6105);
	not 	XG2555 	(g7841,g904);
	not 	XG2556 	(g10078,g1854);
	not 	XG2557 	(g9369,g5084);
	not 	XG2558 	(g9036,g5084);
	not 	XG2559 	(I12890,g4219);
	nor 	XG2560 	(g9762,g2421,g2495);
	not 	XG2561 	(g7456,g2495);
	not 	XG2562 	(g9546,g2437);
	not 	XG2563 	(g10217,g2102);
	not 	XG2564 	(g8205,g2208);
	not 	XG2565 	(g9834,g2579);
	nor 	XG2566 	(g7781,g4057,g4064);
	nand 	XG2567 	(g7611,g4064,g4057);
	not 	XG2568 	(g7927,g4064);
	not 	XG2569 	(g7650,g4064);
	nor 	XG2570 	(g8984,g4975,g4899);
	not 	XG2571 	(g6992,g4899);
	not 	XG2572 	(g8938,g4899);
	not 	XG2573 	(I12183,g2719);
	not 	XG2574 	(g9354,g2719);
	not 	XG2575 	(g8796,g4785);
	not 	XG2576 	(g8774,g781);
	not 	XG2577 	(I12049,g781);
	not 	XG2578 	(g9891,g6173);
	not 	XG2579 	(I16803,g6369);
	and 	XG2580 	(g8583,g2912,g2917);
	not 	XG2581 	(g8680,g686);
	not 	XG2582 	(g7957,g1252);
	not 	XG2583 	(g8858,g671);
	not 	XG2584 	(g9759,g2265);
	not 	XG2585 	(I18835,g6365);
	not 	XG2586 	(g7393,g5320);
	not 	XG2587 	(I18647,g5320);
	not 	XG2588 	(g10172,g6459);
	not 	XG2589 	(g9381,g5527);
	not 	XG2590 	(g10206,g4489);
	not 	XG2591 	(g9827,g1974);
	not 	XG2592 	(g7349,g1270);
	not 	XG2593 	(g7953,g4966);
	not 	XG2594 	(g7345,g6415);
	not 	XG2595 	(g9569,g6227);
	not 	XG2596 	(g9863,g5503);
	or 	XG2597 	(g9984,g4242,g4300);
	not 	XG2598 	(g6956,g4242);
	nand 	XG2599 	(I12251,g1129,g1124);
	not 	XG2600 	(g6996,g4955);
	not 	XG2601 	(g9541,g2012);
	not 	XG2602 	(g9326,g6203);
	nand 	XG2603 	(I13043,g5120,g5115);
	not 	XG2604 	(g7392,g4438);
	not 	XG2605 	(g9416,g2429);
	not 	XG2606 	(g8655,g2787);
	not 	XG2607 	(g10156,g2675);
	not 	XG2608 	(I11980,g66);
	not 	XG2609 	(I13326,g66);
	not 	XG2610 	(g8400,g4836);
	not 	XG2611 	(g7716,g1199);
	not 	XG2612 	(g8506,g3782);
	not 	XG2613 	(g9892,g6428);
	not 	XG2614 	(g10200,g2138);
	or 	XG2615 	(g8957,g2357,g2338);
	not 	XG2616 	(I12896,g4229);
	not 	XG2617 	(g7880,g1291);
	not 	XG2618 	(g9492,g2759);
	not 	XG2619 	(I11809,g6741);
	not 	XG2620 	(g10194,g6741);
	not 	XG2621 	(I12070,g785);
	not 	XG2622 	(g8948,g785);
	not 	XG2623 	(g7487,g1259);
	not 	XG2624 	(g8164,g3484);
	not 	XG2625 	(g9269,g5517);
	not 	XG2626 	(g9833,g2449);
	not 	XG2627 	(g9704,g2575);
	not 	XG2628 	(I13007,g65);
	not 	XG2629 	(I12172,g2715);
	not 	XG2630 	(g9285,g2715);
	not 	XG2631 	(g7909,g936);
	not 	XG2632 	(g9848,g4462);
	not 	XG2633 	(I12151,g604);
	not 	XG2634 	(g9044,g604);
	not 	XG2635 	(g9693,g1886);
	nand 	XG2636 	(g10022,g6466,g6474);
	not 	XG2637 	(g9212,g6466);
	not 	XG2638 	(g9626,g6466);
	not 	XG2639 	(I15717,g6346);
	not 	XG2640 	(g9338,g1870);
	not 	XG2641 	(g10057,g6455);
	not 	XG2642 	(g9014,g3004);
	nand 	XG2643 	(I13390,g1825,g1821);
	not 	XG2644 	(g9824,g1825);
	not 	XG2645 	(g9951,g6133);
	not 	XG2646 	(g7479,g1008);
	not 	XG2647 	(g7178,g4392);
	not 	XG2648 	(I12493,g5002);
	not 	XG2649 	(g8284,g5002);
	not 	XG2650 	(g10085,g1768);
	not 	XG2651 	(g8677,g4854);
	not 	XG2652 	(g9575,g6509);
	not 	XG2653 	(g9690,g732);
	not 	XG2654 	(g6836,g1322);
	nand 	XG2655 	(g9543,g2185,g2217);
	not 	XG2656 	(g8150,g2185);
	not 	XG2657 	(g8607,g37);
	not 	XG2658 	(I17970,g4027);
	nor 	XG2659 	(g9755,g1996,g2070);
	not 	XG2660 	(g7451,g2070);
	not 	XG2661 	(I12463,g4812);
	not 	XG2662 	(g8236,g4812);
	not 	XG2663 	(g9946,g6093);
	not 	XG2664 	(g6837,g968);
	not 	XG2665 	(g7219,g4405);
	not 	XG2666 	(I11892,g4408);
	not 	XG2667 	(g7244,g4408);
	not 	XG2668 	(g9568,g6181);
	not 	XG2669 	(I13539,g6381);
	not 	XG2670 	(g10053,g6381);
	not 	XG2671 	(g6988,g4765);
	not 	XG2672 	(g7943,g1395);
	or 	XG2673 	(g8956,g1932,g1913);
	not 	XG2674 	(g7380,g2331);
	not 	XG2675 	(I12534,g50);
	not 	XG2676 	(g7592,g347);
	not 	XG2677 	(g9501,g5731);
	not 	XG2678 	(I11734,g4473);
	not 	XG2679 	(g7873,g1266);
	not 	XG2680 	(g9443,g5489);
	nand 	XG2681 	(g8769,g714,g691);
	not 	XG2682 	(g6811,g714);
	not 	XG2683 	(g9766,g2748);
	not 	XG2684 	(I12056,g2748);
	not 	XG2685 	(g9380,g5471);
	not 	XG2686 	(g9761,g2445);
	not 	XG2687 	(g9542,g2173);
	nand 	XG2688 	(I12728,g4287,g4291);
	not 	XG2689 	(I12950,g4287);
	not 	XG2690 	(g9020,g4287);
	or 	XG2691 	(g9013,g2491,g2472);
	nand 	XG2692 	(g7701,g4843,g4849,g4859);
	not 	XG2693 	(g7693,g4849);
	not 	XG2694 	(g9415,g2169);
	not 	XG2695 	(g6847,g2283);
	not 	XG2696 	(g10115,g2283);
	not 	XG2697 	(I13552,g121);
	not 	XG2698 	(g10083,g2407);
	not 	XG2699 	(g8195,g1783);
	not 	XG2700 	(I17932,g3310);
	not 	XG2701 	(g9599,g3310);
	or 	XG2702 	(g9536,g1312,g1351);
	not 	XG2703 	(g7922,g1312);
	not 	XG2704 	(I13634,g79);
	not 	XG2705 	(g8807,g79);
	not 	XG2706 	(g7374,g2227);
	not 	XG2707 	(g9890,g6058);
	not 	XG2708 	(I12773,g4204);
	nand 	XG2709 	(I13401,g2250,g2246);
	not 	XG2710 	(g7998,g392);
	not 	XG2711 	(g7252,g1592);
	not 	XG2712 	(g7212,g6411);
	not 	XG2713 	(g9197,g1221);
	not 	XG2714 	(I13672,g106);
	not 	XG2715 	(g8990,g146);
	not 	XG2716 	(g8290,g218);
	not 	XG2717 	(g6826,g218);
	not 	XG2718 	(g9960,g6474);
	not 	XG2719 	(g8093,g1624);
	nand 	XG2720 	(g7150,g5062,g5016);
	not 	XG2721 	(g9613,g5062);
	not 	XG2722 	(g9309,g5462);
	and 	XG2723 	(g7520,g2689,g2697,g2704);
	nor 	XG2724 	(g7142,g6565,g6573);
	not 	XG2725 	(g9631,g6573);
	nand 	XG2726 	(g9645,g2028,g2060);
	not 	XG2727 	(g8255,g2028);
	not 	XG2728 	(g10042,g2671);
	not 	XG2729 	(I12227,g34);
	not 	XG2730 	(g10037,g1848);
	not 	XG2731 	(g6870,g3089);
	not 	XG2732 	(g8219,g3731);
	not 	XG2733 	(g6999,g86);
	not 	XG2734 	(I13329,g86);
	not 	XG2735 	(g9805,g5485);
	not 	XG2736 	(g9708,g2741);
	not 	XG2737 	(I12041,g2741);
	not 	XG2738 	(g7643,g4322);
	not 	XG2739 	(g9920,g4322);
	not 	XG2740 	(I12907,g4322);
	not 	XG2741 	(I12808,g4322);
	not 	XG2742 	(g9910,g2108);
	not 	XG2743 	(g7195,g25);
	not 	XG2744 	(g8808,g595);
	not 	XG2745 	(I12030,g595);
	not 	XG2746 	(g8259,g2217);
	not 	XG2747 	(g6829,g1319);
	not 	XG2748 	(g10289,g1319);
	not 	XG2749 	(g7854,g1152);
	not 	XG2750 	(g7327,g2165);
	not 	XG2751 	(g9598,g2571);
	not 	XG2752 	(I12167,g5176);
	not 	XG2753 	(g9259,g5176);
	not 	XG2754 	(g6801,g391);
	not 	XG2755 	(g8404,g5005);
	not 	XG2756 	(I12568,g5005);
	not 	XG2757 	(g6855,g2711);
	not 	XG2758 	(g8052,g1211);
	not 	XG2759 	(g9621,g6423);
	not 	XG2760 	(g6993,g4859);
	not 	XG2761 	(g8714,g4859);
	not 	XG2762 	(g8181,g424);
	not 	XG2763 	(g7553,g1274);
	not 	XG2764 	(I13740,g85);
	not 	XG2765 	(g8616,g2803);
	not 	XG2766 	(g10059,g6451);
	not 	XG2767 	(g10117,g2509);
	not 	XG2768 	(g9776,g5073);
	not 	XG2769 	(g7939,g1280);
	not 	XG2770 	(g8354,g4815);
	not 	XG2771 	(I12530,g4815);
	not 	XG2772 	(g9299,g5124);
	not 	XG2773 	(g9778,g5069);
	not 	XG2774 	(g9072,g2994);
	not 	XG2775 	(g7891,g2994);
	not 	XG2776 	(g7268,g1636);
	not 	XG2777 	(g9971,g2093);
	not 	XG2778 	(g10213,g6732);
	not 	XG2779 	(g7533,g1306);
	not 	XG2780 	(g7247,g5377);
	not 	XG2781 	(g7936,g1061);
	not 	XG2782 	(g9698,g2181);
	nand 	XG2783 	(I12269,g956,g1141);
	not 	XG2784 	(g6817,g956);
	not 	XG2785 	(g9692,g1756);
	not 	XG2786 	(g9934,g5849);
	not 	XG2787 	(g10204,g2685);
	not 	XG2788 	(g6854,g2685);
	not 	XG2789 	(g7328,g2197);
	nand 	XG2790 	(g9567,g6120,g6116);
	not 	XG2791 	(g9516,g6116);
	not 	XG2792 	(g7387,g2421);
	not 	XG2793 	(g7972,g1046);
	not 	XG2794 	(g6819,g1046);
	not 	XG2795 	(g8183,g482);
	not 	XG2796 	(g9467,g6434);
	not 	XG2797 	(g8466,g1514);
	not 	XG2798 	(g7440,g329);
	not 	XG2799 	(g9576,g6565);
	not 	XG2800 	(g7649,g1345);
	not 	XG2801 	(g9685,g6533);
	not 	XG2802 	(g9842,g3274);
	not 	XG2803 	(I17814,g3274);
	not 	XG2804 	(g8431,g3085);
	not 	XG2805 	(g7888,g1536);
	not 	XG2806 	(g8944,g370);
	not 	XG2807 	(g10130,g5694);
	not 	XG2808 	(g10111,g1858);
	not 	XG2809 	(g6839,g1858);
	not 	XG2810 	(g6998,g4932);
	not 	XG2811 	(g8440,g3431);
	not 	XG2812 	(g8064,g3376);
	not 	XG2813 	(g9653,g2441);
	not 	XG2814 	(g7361,g1874);
	and 	XG2815 	(g10290,g4349,g4358);
	not 	XG2816 	(g8977,g4349);
	not 	XG2817 	(I12930,g4349);
	not 	XG2818 	(I12826,g4349);
	not 	XG2819 	(g7992,g5008);
	not 	XG2820 	(g9909,g1978);
	not 	XG2821 	(g9484,g1612);
	not 	XG2822 	(I13057,g112);
	not 	XG2823 	(g10019,g6479);
	not 	XG2824 	(g10080,g1982);
	not 	XG2825 	(I18667,g6661);
	not 	XG2826 	(g7522,g6661);
	not 	XG2827 	(g10212,g6390);
	not 	XG2828 	(g7752,g1542);
	not 	XG2829 	(g8872,g4258);
	not 	XG2830 	(g8514,g4258);
	not 	XG2831 	(g7971,g4818);
	not 	XG2832 	(g7239,g5033);
	not 	XG2833 	(g8088,g1554);
	not 	XG2834 	(g8594,g3849);
	not 	XG2835 	(g7514,g6704);
	not 	XG2836 	(I18778,g6704);
	not 	XG2837 	(g7050,g5845);
	not 	XG2838 	(g9619,g5845);
	not 	XG2839 	(g8822,g4975);
	not 	XG2840 	(I12092,g790);
	not 	XG2841 	(g9003,g790);
	not 	XG2842 	(g10120,g1902);
	not 	XG2843 	(g9517,g6163);
	not 	XG2844 	(g7835,g4125);
	not 	XG2845 	(g7040,g4821);
	not 	XG2846 	(g8741,g4821);
	not 	XG2847 	(g8676,g4821);
	not 	XG2848 	(g10335,g4483);
	not 	XG2849 	(g9373,g5142);
	not 	XG2850 	(g10178,g2126);
	not 	XG2851 	(g6845,g2126);
	not 	XG2852 	(g8697,g3694);
	not 	XG2853 	(g9732,g5481);
	not 	XG2854 	(g9721,g5097);
	not 	XG2855 	(I11843,g111);
	not 	XG2856 	(g7222,g4427);
	not 	XG2857 	(g9963,g7);
	nand 	XG2858 	(I12876,g4180,g4200);
	not 	XG2859 	(I12770,g4200);
	not 	XG2860 	(g10035,g1720);
	not 	XG2861 	(g7534,g1367);
	not 	XG2862 	(g9777,g5112);
	not 	XG2863 	(I11629,g19);
	not 	XG2864 	(g10140,g19);
	not 	XG2865 	(I11721,g4145);
	not 	XG2866 	(g9284,g2161);
	not 	XG2867 	(g8890,g376);
	not 	XG2868 	(g7418,g2361);
	not 	XG2869 	(I12000,g582);
	not 	XG2870 	(g8891,g582);
	not 	XG2871 	(g8310,g2051);
	not 	XG2872 	(g7870,g1193);
	not 	XG2873 	(g9792,g5401);
	not 	XG2874 	(g8540,g3408);
	not 	XG2875 	(g10121,g2327);
	not 	XG2876 	(g7933,g907);
	not 	XG2877 	(g7858,g947);
	not 	XG2878 	(g10177,g1834);
	not 	XG2879 	(g9386,g5727);
	not 	XG2880 	(g9489,g2303);
	not 	XG2881 	(g8620,g3065);
	not 	XG2882 	(g6810,g723);
	not 	XG2883 	(g9282,g723);
	not 	XG2884 	(I11785,g5703);
	not 	XG2885 	(g10093,g5703);
	not 	XG2886 	(g10014,g6439);
	not 	XG2887 	(g7314,g1740);
	not 	XG2888 	(g8346,g3845);
	not 	XG2889 	(g6927,g3845);
	not 	XG2890 	(g10114,g2116);
	nand 	XG2891 	(I13334,g1691,g1687);
	not 	XG2892 	(g10182,g2681);
	not 	XG2893 	(g9914,g2533);
	not 	XG2894 	(g7802,g324);
	not 	XG2895 	(g10219,g2697);
	not 	XG2896 	(g9875,g5747);
	not 	XG2897 	(I13597,g4417);
	not 	XG2898 	(I12214,g6561);
	not 	XG2899 	(g9529,g6561);
	not 	XG2900 	(g10116,g2413);
	not 	XG2901 	(g9751,g1710);
	not 	XG2902 	(g9630,g6527);
	not 	XG2903 	(g9961,g6404);
	not 	XG2904 	(g9749,g1691);
	not 	XG2905 	(g9924,g5644);
	not 	XG2906 	(g7041,g5644);
	not 	XG2907 	(g7003,g5152);
	not 	XG2908 	(g9499,g5152);
	not 	XG2909 	(g10129,g5352);
	not 	XG2910 	(g9564,g6120);
	not 	XG2911 	(g9184,g6120);
	not 	XG2912 	(g8612,g2775);
	not 	XG2913 	(I17787,g3267);
	not 	XG2914 	(g9660,g3267);
	not 	XG2915 	(g8365,g2060);
	not 	XG2916 	(g8396,g3401);
	not 	XG2917 	(g7805,g4366);
	not 	XG2918 	(I13548,g94);
	not 	XG2919 	(g8439,g3129);
	not 	XG2920 	(I17892,g3325);
	not 	XG2921 	(g9234,g5170);
	not 	XG2922 	(g9740,g5821);
	not 	XG2923 	(g8119,g3727);
	not 	XG2924 	(g6983,g4698);
	not 	XG2925 	(g8666,g3703);
	not 	XG2926 	(I11708,g3703);
	not 	XG2927 	(g9247,g1559);
	not 	XG2928 	(g8137,g411);
	not 	XG2929 	(g8057,g3068);
	not 	XG2930 	(g6850,g2704);
	not 	XG2931 	(g9995,g6035);
	not 	XG2932 	(I13483,g6035);
	not 	XG2933 	(g9809,g6082);
	not 	XG2934 	(I12497,g49);
	not 	XG2935 	(g6828,g1300);
	not 	XG2936 	(g8451,g4057);
	not 	XG2937 	(g8630,g4843);
	not 	XG2938 	(g9607,g5046);
	not 	XG2939 	(g9829,g2250);
	not 	XG2940 	(g8273,g2453);
	not 	XG2941 	(g9558,g5841);
	not 	XG2942 	(g9931,g5763);
	not 	XG2943 	(g8553,g3747);
	not 	XG2944 	(g9037,g164);
	not 	XG2945 	(I12128,g4253);
	not 	XG2946 	(g10337,g5016);
	not 	XG2947 	(g8341,g3119);
	not 	XG2948 	(g7503,g1351);
	not 	XG2949 	(g8139,g1648);
	not 	XG2950 	(I11740,g4519);
	not 	XG2951 	(g9257,g5115);
	not 	XG2952 	(I11697,g3352);
	not 	XG2953 	(g8644,g3352);
	not 	XG2954 	(g6815,g929);
	not 	XG2955 	(g8389,g3125);
	not 	XG2956 	(g8450,g3821);
	not 	XG2957 	(g8509,g4141);
	not 	XG2958 	(I11746,g4570);
	not 	XG2959 	(g9547,g2735);
	not 	XG2960 	(g10147,g728);
	not 	XG2961 	(g9860,g5417);
	not 	XG2962 	(g10231,g2661);
	not 	XG2963 	(g10112,g1988);
	not 	XG2964 	(g9614,g5128);
	not 	XG2965 	(g9200,g1548);
	not 	XG2966 	(g8009,g3106);
	not 	XG2967 	(g7686,g4659);
	not 	XG2968 	(g9024,g4358);
	not 	XG2969 	(I12954,g4358);
	not 	XG2970 	(g8241,g1792);
	not 	XG2971 	(g10113,g2084);
	not 	XG2972 	(g8477,g3061);
	not 	XG2973 	(I12855,g4311);
	not 	XG2974 	(g7166,g4311);
	not 	XG2975 	(g7627,g4311);
	not 	XG2976 	(I12823,g4311);
	not 	XG2977 	(g9843,g4311);
	not 	XG2978 	(I12787,g4311);
	not 	XG2979 	(g9915,g2583);
	not 	XG2980 	(g8282,g3841);
	not 	XG2981 	(I12709,g4284);
	not 	XG2982 	(g8591,g3763);
	not 	XG2983 	(g9983,g4239);
	not 	XG2984 	(g8016,g3391);
	not 	XG2985 	(g8912,g4180);
	not 	XG2986 	(g8744,g691);
	not 	XG2987 	(g9731,g5366);
	not 	XG2988 	(g8993,g385);
	not 	XG2989 	(g9414,g2004);
	not 	XG2990 	(g10218,g2527);
	not 	XG2991 	(g9804,g5456);
	not 	XG2992 	(g6959,g4420);
	not 	XG2993 	(g10334,g4420);
	not 	XG2994 	(g9433,g5148);
	not 	XG2995 	(g6975,g4507);
	not 	XG2996 	(g10090,g5348);
	not 	XG2997 	(g10165,g5698);
	not 	XG2998 	(g8647,g3416);
	not 	XG2999 	(g7751,g1521);
	not 	XG3000 	(g8114,g3522);
	not 	XG3001 	(g8058,g3115);
	not 	XG3002 	(I11617,g1);
	not 	XG3003 	(I11620,g1);
	not 	XG3004 	(g6960,g1);
	not 	XG3005 	(g10278,g4628);
	not 	XG3006 	(g7369,g1996);
	not 	XG3007 	(g8130,g4515);
	not 	XG3008 	(g10077,g1724);
	not 	XG3009 	(g6838,g1724);
	not 	XG3010 	(g7581,g1379);
	not 	XG3011 	(I12987,g12);
	not 	XG3012 	(g7115,g12);
	not 	XG3013 	(g9488,g1878);
	not 	XG3014 	(I13715,g71);
	not 	XG3015 	(I12799,g59);
	not 	XG3016 	(I12712,g59);
	not 	XG3017 	(g10430,I13847);
	not 	XG3018 	(g10364,g6869);
	not 	XG3019 	(g12076,g9280);
	not 	XG3020 	(g12180,g9477);
	not 	XG3021 	(g12181,g9478);
	not 	XG3022 	(g12036,g9245);
	not 	XG3023 	(g11964,g9154);
	not 	XG3024 	(g11984,g9186);
	not 	XG3025 	(g12012,g9213);
	not 	XG3026 	(g12321,g9637);
	not 	XG3027 	(g11963,g9153);
	not 	XG3028 	(g11912,g8989);
	not 	XG3029 	(g12074,I14932);
	not 	XG3030 	(g12217,I15070);
	not 	XG3031 	(g10877,I14079);
	not 	XG3032 	(g11988,I14836);
	not 	XG3033 	(g12109,I14967);
	not 	XG3034 	(g12038,I14896);
	not 	XG3035 	(g11165,I14222);
	not 	XG3036 	(g12143,I14999);
	not 	XG3037 	(g12037,I14893);
	not 	XG3038 	(g11204,I14271);
	not 	XG3039 	(g11949,I14773);
	not 	XG3040 	(g12322,I15162);
	not 	XG3041 	(g11235,I14301);
	not 	XG3042 	(g12075,I14935);
	not 	XG3043 	(g11182,I14241);
	not 	XG3044 	(g11989,I14839);
	not 	XG3045 	(g12041,I14905);
	not 	XG3046 	(g12013,I14866);
	not 	XG3047 	(g12182,I15030);
	not 	XG3048 	(g11965,I14797);
	not 	XG3049 	(g12040,I14902);
	not 	XG3050 	(g12218,I15073);
	not 	XG3051 	(g11928,I14742);
	not 	XG3052 	(g12110,I14970);
	not 	XG3053 	(g11867,I14679);
	not 	XG3054 	(g11985,I14827);
	not 	XG3055 	(g8712,I12712);
	not 	XG3056 	(g8805,I12799);
	not 	XG3057 	(g10287,I13715);
	nand 	XG3058 	(g10520,g7115,g7195);
	not 	XG3059 	(g9104,I12987);
	nor 	XG3060 	(g11869,g7581,g7534,g7649);
	nand 	XG3061 	(g10603,g9751,g10077);
	nand 	XG3062 	(g10585,g7451,g1996);
	not 	XG3063 	(g10380,g6960);
	not 	XG3064 	(g6755,I11620);
	not 	XG3065 	(g6754,I11617);
	nor 	XG3066 	(g11618,g8070,g8114);
	nor 	XG3067 	(g11527,g8114,g8165);
	nor 	XG3068 	(g11483,g3522,g8165);
	and 	XG3069 	(g12220,g7535,g1521);
	nand 	XG3070 	(g12294,g10090,g7018,g10044);
	nand 	XG3071 	(I15128,g2527,g9914);
	nand 	XG3072 	(I14609,g8678,g8993);
	nand 	XG3073 	(g10537,g5366,g7138);
	not 	XG3074 	(I13995,g8744);
	not 	XG3075 	(I14033,g8912);
	nand 	XG3076 	(I12878,I12876,g4180);
	nor 	XG3077 	(g11414,g8593,g8591);
	nor 	XG3078 	(g11360,g8669,g3763);
	not 	XG3079 	(g8703,I12709);
	nand 	XG3080 	(I12204,I12203,g1094);
	not 	XG3081 	(g8791,I12787);
	nand 	XG3082 	(g10820,g9843,g9920,g9985);
	not 	XG3083 	(g8841,I12823);
	nand 	XG3084 	(g12797,g7627,g7643,g7655,g10275);
	and 	XG3085 	(g11018,g7627,g7643,g7655);
	not 	XG3086 	(g8876,I12855);
	nor 	XG3087 	(g11345,g8479,g8477);
	nor 	XG3088 	(g11273,g8620,g3061);
	nor 	XG3089 	(g12117,g9755,g10113);
	nand 	XG3090 	(g12114,g8146,g8241);
	nand 	XG3091 	(g11953,g8241,g8195);
	nand 	XG3092 	(g12079,g8195,g1792);
	not 	XG3093 	(g9021,I12954);
	nand 	XG3094 	(g10614,g8928,g8977,g9024);
	and 	XG3095 	(g12687,g8977,g9024);
	and 	XG3096 	(g12762,g8977,g4358);
	nor 	XG3097 	(g11006,g7836,g7686);
	nand 	XG3098 	(I12345,I12344,g3106);
	nor 	XG3099 	(g11171,g9091,g9200,g9226,g8088);
	and 	XG3100 	(g10921,g8685,g1548);
	nand 	XG3101 	(I14712,g5128,g9671);
	nand 	XG3102 	(I15174,g2661,g9977);
	nor 	XG3103 	(g12296,g9862,g9860);
	nor 	XG3104 	(g12201,g10047,g5417);
	nand 	XG3105 	(g11708,g10110,g10147);
	not 	XG3106 	(g6974,I11746);
	nor 	XG3107 	(g10808,g7611,g8509);
	and 	XG3108 	(g10998,g7650,g8451,g8509,g8567);
	and 	XG3109 	(g10841,g8567,g8509);
	and 	XG3110 	(g10677,g7611,g4141);
	nand 	XG3111 	(I14204,g3821,g8508);
	nand 	XG3112 	(g11382,g8663,g6895,g8644);
	not 	XG3113 	(g6875,I11697);
	nand 	XG3114 	(I13044,I13043,g5115);
	not 	XG3115 	(g6972,I11740);
	nand 	XG3116 	(g11934,g8187,g8139);
	nand 	XG3117 	(g12016,g8093,g1648);
	nand 	XG3118 	(g11914,g1648,g8187);
	nor 	XG3119 	(g12113,g8187,g1648);
	and 	XG3120 	(g12817,g7601,g1351);
	and 	XG3121 	(g11366,g10338,g5016);
	not 	XG3122 	(g7640,I12128);
	and 	XG3123 	(I24033,g3747,g8443,g8219);
	and 	XG3124 	(I24054,g3747,g8075,g8443);
	nor 	XG3125 	(g12346,g9933,g9931);
	nor 	XG3126 	(g12249,g10096,g5763);
	nand 	XG3127 	(g12194,g8273,g8373);
	nand 	XG3128 	(g12225,g2453,g8324);
	nand 	XG3129 	(g12023,g8373,g2453);
	nor 	XG3130 	(g12483,g8324,g2453);
	nand 	XG3131 	(I13403,I13401,g2250);
	nor 	XG3132 	(g10884,g8451,g7650);
	and 	XG3133 	(g10626,g7927,g4057);
	nor 	XG3134 	(g10922,g4057,g7650);
	and 	XG3135 	(g11003,g1300,g7880);
	nand 	XG3136 	(I12289,I12287,g1300);
	not 	XG3137 	(g8285,I12497);
	not 	XG3138 	(g9935,I13483);
	nor 	XG3139 	(g12252,g10185,g9995);
	not 	XG3140 	(g12830,g9995);
	and 	XG3141 	(g11126,g10185,g6035);
	not 	XG3142 	(g10362,g6850);
	and 	XG3143 	(g10684,g411,g7998);
	not 	XG3144 	(g6905,I11708);
	nand 	XG3145 	(g11412,g8697,g6918,g8666);
	not 	XG3146 	(g10388,g6983);
	and 	XG3147 	(g11010,g8933,g4698);
	nand 	XG3148 	(g12292,g8933,g4698);
	nand 	XG3149 	(I14764,g5821,g9808);
	nor 	XG3150 	(g12235,g9206,g9234);
	nor 	XG3151 	(g12646,g9206,g9234);
	nor 	XG3152 	(g12553,g9206,g5170);
	and 	XG3153 	(g11205,g8439,g8217);
	not 	XG3154 	(g10029,I13548);
	nand 	XG3155 	(g12190,g8255,g8365);
	nand 	XG3156 	(g11994,g8365,g8310);
	nand 	XG3157 	(g12148,g8310,g2060);
	nand 	XG3158 	(g11441,g3267,g9599);
	nand 	XG3159 	(I12241,I12240,g1111);
	and 	XG3160 	(g11046,g6120,g9889);
	and 	XG3161 	(g12027,g9729,g9499);
	nand 	XG3162 	(g12344,g10130,g7041,g10093);
	not 	XG3163 	(g10401,g7041);
	nand 	XG3164 	(I13336,I13334,g1691);
	nand 	XG3165 	(g10598,g6404,g7191);
	nand 	XG3166 	(I14991,g6527,g9685);
	nand 	XG3167 	(I12270,I12269,g1141);
	nor 	XG3168 	(g12752,g9529,g9576);
	not 	XG3169 	(g10581,g9529);
	not 	XG3170 	(g7812,I12214);
	not 	XG3171 	(g10087,I13597);
	and 	XG3172 	(I24530,g5747,g9733,g9501);
	and 	XG3173 	(I24552,g5747,g9316,g9733);
	nand 	XG3174 	(g10759,g324,g7537);
	nand 	XG3175 	(I15333,g2116,g10152);
	and 	XG3176 	(g11244,g8566,g8346);
	nor 	XG3177 	(g11954,g7314,g9538);
	and 	XG3178 	(I24603,g6439,g9467,g9892);
	and 	XG3179 	(I24585,g6439,g9892,g9621);
	not 	XG3180 	(g7028,I11785);
	nand 	XG3181 	(I15041,g1834,g9752);
	nor 	XG3182 	(g11384,g8540,g8538);
	and 	XG3183 	(I24508,g5401,g9672,g9434);
	and 	XG3184 	(I24527,g5401,g9264,g9672);
	nand 	XG3185 	(g11330,g1193,g9483);
	nand 	XG3186 	(g12116,g8255,g2051);
	not 	XG3187 	(g7515,I12000);
	nand 	XG3188 	(g10586,g7418,g7380);
	and 	XG3189 	(g11939,g7380,g2361);
	nand 	XG3190 	(I14350,g8848,g8890);
	nor 	XG3191 	(g11607,g376,g8993,g8848);
	not 	XG3192 	(g6946,I11721);
	not 	XG3193 	(I14505,g10140);
	not 	XG3194 	(g6772,I11629);
	nand 	XG3195 	(I12877,I12876,g4200);
	not 	XG3196 	(I14050,g9963);
	not 	XG3197 	(g7161,I11843);
	nor 	XG3198 	(g12160,g9724,g9721);
	and 	XG3199 	(g11027,g9724,g5097);
	nand 	XG3200 	(g10622,g9973,g10178);
	nor 	XG3201 	(g12228,g10335,g10184,g10206,g10222);
	not 	XG3202 	(g10403,g7040);
	not 	XG3203 	(I14267,g7835);
	nor 	XG3204 	(g11201,g7765,g4125);
	not 	XG3205 	(g7618,I12092);
	nor 	XG3206 	(g11834,g8822,g8938);
	nor 	XG3207 	(g11804,g4975,g8938);
	and 	XG3208 	(g12099,g9888,g9619);
	nand 	XG3209 	(g12476,g6704,g7498);
	nand 	XG3210 	(g10556,g8133,g7971);
	and 	XG3211 	(g10827,g4258,g8914);
	nor 	XG3212 	(g12358,g10022,g10019);
	and 	XG3213 	(g11127,g10022,g6479);
	not 	XG3214 	(g9281,I13057);
	nand 	XG3215 	(g10617,g9909,g10151);
	nand 	XG3216 	(g10573,g8179,g7992);
	not 	XG3217 	(g8844,I12826);
	not 	XG3218 	(g8974,I12930);
	nor 	XG3219 	(g11972,g7361,g9591);
	and 	XG3220 	(g10625,g7926,g3431);
	nand 	XG3221 	(g10609,g9826,g10111);
	nand 	XG3222 	(I14508,g8721,g370);
	nand 	XG3223 	(g11374,g1536,g9536);
	nor 	XG3224 	(g11270,g8434,g8431);
	and 	XG3225 	(g10654,g8434,g3085);
	and 	XG3226 	(g12043,g7601,g1345);
	nor 	XG3227 	(g12680,g9576,g9631);
	nor 	XG3228 	(g12632,g6565,g9631);
	nor 	XG3229 	(g10715,g8466,g8526);
	nor 	XG3230 	(g10699,g1514,g8526);
	nand 	XG3231 	(I11866,I11864,g4401);
	not 	XG3232 	(g10356,g6819);
	nor 	XG3233 	(g10760,g7479,g1046);
	nand 	XG3234 	(g10587,g7456,g2421);
	nand 	XG3235 	(g10568,g7374,g7328);
	nand 	XG3236 	(g11996,g2197,g7280);
	nand 	XG3237 	(g10653,g10042,g10204);
	nand 	XG3238 	(I12271,I12269,g956);
	nand 	XG3239 	(I12374,I12372,g3462);
	nand 	XG3240 	(g12526,g10213,g7110,g10194);
	nand 	XG3241 	(I13511,I13509,g2093);
	nand 	XG3242 	(g10550,g7308,g7268);
	nand 	XG3243 	(g11969,g1636,g7252);
	nor 	XG3244 	(g10615,g7308,g1636);
	nor 	XG3245 	(g12234,g9778,g9776);
	nor 	XG3246 	(g12126,g5069,g9989);
	nor 	XG3247 	(g12163,g9989,g5073);
	nor 	XG3248 	(g12121,g9762,g10117);
	nand 	XG3249 	(I13391,I13390,g1821);
	nor 	XG3250 	(g12466,g10059,g10057);
	nor 	XG3251 	(g12318,g6451,g10172);
	not 	XG3252 	(g10319,I13740);
	and 	XG3253 	(g10565,g424,g8182);
	nor 	XG3254 	(g11148,g9050,g9174,g9197,g8052);
	nor 	XG3255 	(g12550,g9259,g9300);
	not 	XG3256 	(g10489,g9259);
	not 	XG3257 	(g7704,I12167);
	nor 	XG3258 	(g11958,g7327,g9543);
	not 	XG3259 	(g11017,g10289);
	nand 	XG3260 	(g11957,g8259,g8205);
	nand 	XG3261 	(g12118,g8150,g8259);
	nand 	XG3262 	(g12083,g8205,g2217);
	not 	XG3263 	(g7542,I12030);
	not 	XG3264 	(g8818,I12808);
	not 	XG3265 	(g8922,I12907);
	not 	XG3266 	(g12399,g9920);
	not 	XG3267 	(g7558,I12041);
	nand 	XG3268 	(g12289,g9708,g9766,g9978);
	not 	XG3269 	(I14567,g9708);
	and 	XG3270 	(g12065,g9805,g9557);
	not 	XG3271 	(g9747,I13329);
	not 	XG3272 	(g10398,g6999);
	not 	XG3273 	(g10367,g6870);
	nand 	XG3274 	(I15253,g1848,g10078);
	not 	XG3275 	(g7831,I12227);
	nor 	XG3276 	(g11995,g7410,g9645);
	not 	XG3277 	(g12082,g9645);
	not 	XG3278 	(g10428,g9631);
	nand 	XG3279 	(I13078,I13077,g5462);
	nor 	XG3280 	(g11862,g7150,g7134);
	nand 	XG3281 	(g12078,g8093,g8187);
	nand 	XG3282 	(g11952,g8187,g1624);
	and 	XG3283 	(g11047,g9212,g6474);
	not 	XG3284 	(g10198,I13672);
	and 	XG3285 	(g10934,g7918,g9197);
	nand 	XG3286 	(g11130,g7918,g1221);
	nor 	XG3287 	(g11945,g7228,g7212);
	nand 	XG3288 	(I13184,I13182,g6505);
	nand 	XG3289 	(g10529,g7308,g1592);
	nor 	XG3290 	(g11216,g8037,g7998);
	nand 	XG3291 	(I12470,I12468,g392);
	nand 	XG3292 	(g10578,g6058,g7174);
	nand 	XG3293 	(I12253,I12251,g1129);
	not 	XG3294 	(g10141,I13634);
	nand 	XG3295 	(I12729,I12728,g4291);
	nor 	XG3296 	(g11469,g645,g9903,g650);
	and 	XG3297 	(g12795,g7601,g1312);
	nand 	XG3298 	(g11355,g3310,g9551);
	nand 	XG3299 	(g12045,g8146,g1783);
	not 	XG3300 	(g10031,I13552);
	nand 	XG3301 	(g10611,g9831,g10115);
	nor 	XG3302 	(g11012,g7846,g7693);
	nor 	XG3303 	(g10862,g7840,g7701);
	not 	XG3304 	(g12088,g7701);
	nor 	XG3305 	(g12486,g8905,g8957,g9013,g9055);
	nand 	XG3306 	(I12730,I12728,g4287);
	not 	XG3307 	(g7586,I12056);
	not 	XG3308 	(I14584,g9766);
	not 	XG3309 	(g10354,g6811);
	nand 	XG3310 	(I14883,g5489,g9500);
	not 	XG3311 	(g6961,I11734);
	nor 	XG3312 	(g10799,g7541,g347);
	not 	XG3313 	(g8355,I12534);
	nand 	XG3314 	(g12022,g2331,g7335);
	nor 	XG3315 	(g12435,g8863,g8904,g8956,g9012);
	not 	XG3316 	(g10391,g6988);
	nor 	XG3317 	(g12314,g10207,g10053);
	not 	XG3318 	(g10427,g10053);
	not 	XG3319 	(g10003,I13539);
	and 	XG3320 	(g11142,g10207,g6381);
	nand 	XG3321 	(I14955,g6181,g9620);
	and 	XG3322 	(I13862,g7258,g7219,g7232);
	and 	XG3323 	(I24582,g6093,g9397,g9809);
	and 	XG3324 	(I24555,g6093,g9809,g9559);
	nand 	XG3325 	(g10602,g7451,g7411);
	and 	XG3326 	(g11956,g7411,g2070);
	not 	XG3327 	(I14326,g8607);
	nand 	XG3328 	(g12149,g2185,g8205);
	not 	XG3329 	(g12021,g9543);
	nor 	XG3330 	(g12374,g8205,g2185);
	not 	XG3331 	(g10360,g6836);
	nand 	XG3332 	(I14247,g8091,g1322);
	nand 	XG3333 	(I12098,I12096,g1322);
	and 	XG3334 	(g12794,g7567,g1008);
	nor 	XG3335 	(g12308,g9954,g9951);
	and 	XG3336 	(g11115,g9954,g6133);
	and 	XG3337 	(g10873,g9015,g3004);
	nor 	XG3338 	(g12361,g10172,g6455);
	nand 	XG3339 	(g12523,g6346,g7563);
	not 	XG3340 	(g11911,g10022);
	not 	XG3341 	(g7674,I12151);
	not 	XG3342 	(g7717,I12172);
	not 	XG3343 	(g9185,I13007);
	nor 	XG3344 	(g12695,g9239,g9269);
	nor 	XG3345 	(g12297,g9239,g9269);
	nor 	XG3346 	(g12604,g9239,g5517);
	and 	XG3347 	(g10665,g8292,g209);
	nand 	XG3348 	(I14275,g3484,g8218);
	not 	XG3349 	(g7596,I12070);
	not 	XG3350 	(g7097,I11809);
	and 	XG3351 	(g10656,g7952,g3782);
	not 	XG3352 	(g9746,I13326);
	not 	XG3353 	(g7474,I11980);
	and 	XG3354 	(g10683,g4438,g7289);
	nor 	XG3355 	(g12419,g9326,g9402);
	nor 	XG3356 	(g12780,g9326,g9402);
	not 	XG3357 	(g10519,g9326);
	nor 	XG3358 	(g12744,g6203,g9402);
	not 	XG3359 	(g10387,g6996);
	nand 	XG3360 	(I12252,I12251,g1124);
	not 	XG3361 	(g10349,g6956);
	nor 	XG3362 	(g12622,g9518,g9569);
	not 	XG3363 	(g12831,g9569);
	nor 	XG3364 	(g10421,g9518,g6227);
	nand 	XG3365 	(g11173,g9064,g7898,g4966);
	nor 	XG3366 	(g11232,g9064,g7898,g4966);
	nor 	XG3367 	(g12601,g9311,g9381);
	nor 	XG3368 	(g12505,g9381,g9444);
	nor 	XG3369 	(g12453,g5527,g9444);
	nand 	XG3370 	(g12244,g5320,g7343);
	or 	XG3371 	(g11380,g8530,g8583);
	not 	XG3372 	(g7566,I12049);
	nor 	XG3373 	(g11797,g8796,g8883);
	nor 	XG3374 	(g11773,g4785,g8883);
	not 	XG3375 	(g7753,I12183);
	not 	XG3376 	(g11034,g7611);
	nand 	XG3377 	(g10604,g7456,g7424);
	and 	XG3378 	(g11960,g7424,g2495);
	and 	XG3379 	(g11023,g5084,g9669);
	nor 	XG3380 	(g12418,g10001,g9999);
	nor 	XG3381 	(g12256,g6105,g10136);
	not 	XG3382 	(g10413,g7110);
	not 	XG3383 	(g7595,I12067);
	not 	XG3384 	(g7659,I12141);
	nor 	XG3385 	(g11950,g9166,g9220);
	nor 	XG3386 	(g11913,g9166,g7197);
	nand 	XG3387 	(g11968,g9086,g9334,g837);
	nand 	XG3388 	(g11933,g7197,g9334,g837);
	and 	XG3389 	(g11029,g9103,g5782);
	not 	XG3390 	(I15382,g9071);
	not 	XG3391 	(g7647,I12132);
	not 	XG3392 	(g10377,g6940);
	not 	XG3393 	(g10664,g8928);
	not 	XG3394 	(g8821,I12811);
	not 	XG3395 	(g8879,I12858);
	not 	XG3396 	(g8925,I12910);
	not 	XG3397 	(g8792,I12790);
	and 	XG3398 	(g11449,g7175,g6052);
	nand 	XG3399 	(g12461,g6000,g7536);
	nor 	XG3400 	(g11283,g9064,g4991,g7953);
	nor 	XG3401 	(g11203,g9064,g4991,g4966);
	not 	XG3402 	(g7004,I11777);
	not 	XG3403 	(g9417,I13124);
	not 	XG3404 	(g7624,I12106);
	nor 	XG3405 	(g11940,g10084,g2712);
	nand 	XG3406 	(I12545,I12544,g191);
	nor 	XG3407 	(g11924,g7209,g7187);
	not 	XG3408 	(g12417,g7175);
	nand 	XG3409 	(I15262,g2273,g10081);
	not 	XG3410 	(g7051,I11793);
	nand 	XG3411 	(g12416,g10166,g7064,g10133);
	nand 	XG3412 	(I13453,I13452,g1955);
	not 	XG3413 	(g8085,I12382);
	not 	XG3414 	(g8515,I12631);
	not 	XG3415 	(I14381,g8300);
	and 	XG3416 	(g10624,g3072,g8387);
	nand 	XG3417 	(g10623,g9976,g10181);
	nand 	XG3418 	(g10971,g7886,g7867);
	nand 	XG3419 	(g10946,g7876,g1489);
	nor 	XG3420 	(g12311,g10136,g6109);
	nor 	XG3421 	(g12154,g9835,g10155);
	nand 	XG3422 	(g11172,g3096,g8478);
	not 	XG3423 	(g7565,I12046);
	nand 	XG3424 	(g11279,g3443,g8504);
	nor 	XG3425 	(g12821,g10261,g7149,g10223,g7132);
	nand 	XG3426 	(g12822,g7163,g7224,g7236,g6978);
	not 	XG3427 	(g10383,g6978);
	nor 	XG3428 	(g12364,g10224,g10102);
	not 	XG3429 	(g11948,g10224);
	nand 	XG3430 	(g11881,g3361,g9060);
	not 	XG3431 	(g11383,g9061);
	nand 	XG3432 	(I13464,I13462,g2384);
	nor 	XG3433 	(g11653,g7964,g7980);
	nor 	XG3434 	(g11346,g7964,g7980);
	nor 	XG3435 	(g11566,g7964,g3161);
	nor 	XG3436 	(g11303,g8500,g8497);
	not 	XG3437 	(g11033,g8500);
	nand 	XG3438 	(g10601,g7397,g896);
	not 	XG3439 	(I14158,g8806);
	not 	XG3440 	(g10272,I13705);
	nor 	XG3441 	(g12085,g9700,g10082);
	nor 	XG3442 	(g11935,g7267,g9485);
	not 	XG3443 	(g11991,g9485);
	nand 	XG3444 	(g11998,g8373,g8324);
	nand 	XG3445 	(g11977,g2476,g8373);
	nor 	XG3446 	(g12226,g8373,g2476);
	not 	XG3447 	(g6756,I11623);
	not 	XG3448 	(I14475,g10175);
	not 	XG3449 	(g7543,I12033);
	nor 	XG3450 	(g11846,g7548,g7518,g7635);
	and 	XG3451 	(g12015,g7567,g1002);
	nor 	XG3452 	(g12170,g5413,g10047);
	nand 	XG3453 	(g11020,g9040,g9187);
	nor 	XG3454 	(g11715,g8026,g8080);
	nor 	XG3455 	(g11415,g8026,g8080);
	not 	XG3456 	(g11833,g8026);
	nor 	XG3457 	(g11697,g3857,g8080);
	and 	XG3458 	(g11223,g8505,g8281);
	not 	XG3459 	(g11026,g8434);
	nand 	XG3460 	(I12219,I12217,g1478);
	nand 	XG3461 	(I13498,I13497,g255);
	nor 	XG3462 	(g12050,g9649,g10038);
	nand 	XG3463 	(I15340,g2541,g10154);
	not 	XG3464 	(g10379,g6953);
	not 	XG3465 	(g9917,I13473);
	nor 	XG3466 	(g11107,g9177,g9095);
	not 	XG3467 	(I14054,g10028);
	nand 	XG3468 	(g10796,g7523,g7537);
	nand 	XG3469 	(g10584,g7405,g7362);
	nand 	XG3470 	(g12019,g1906,g7322);
	not 	XG3471 	(g10355,g6816);
	nand 	XG3472 	(I14816,g6513,g9962);
	not 	XG3473 	(g10358,g6827);
	not 	XG3474 	(g7594,I12064);
	not 	XG3475 	(g10582,g7116);
	not 	XG3476 	(g10416,g10318);
	not 	XG3477 	(g9340,I13094);
	not 	XG3478 	(g7117,I11816);
	nand 	XG3479 	(g10755,g1404,g1322,g7675,g7352);
	nand 	XG3480 	(g12415,g5976,g7496);
	not 	XG3481 	(g10288,I13718);
	and 	XG3482 	(g10632,g890,g7441,g7475);
	nor 	XG3483 	(g12739,g9274,g9321);
	nor 	XG3484 	(g12347,g9274,g9321);
	not 	XG3485 	(g10490,g9274);
	nor 	XG3486 	(g12700,g5857,g9321);
	not 	XG3487 	(g12465,g7192);
	not 	XG3488 	(g7615,I12083);
	nor 	XG3489 	(g12025,g7461,g9705);
	nand 	XG3490 	(I13520,I13518,g2518);
	not 	XG3491 	(g10233,I13699);
	nand 	XG3492 	(I12288,I12287,g1484);
	and 	XG3493 	(g10970,g9582,g854);
	nand 	XG3494 	(I11826,I11824,g4601);
	and 	XG3495 	(g12179,g10027,g9745);
	not 	XG3496 	(g10415,g7109);
	nand 	XG3497 	(g10605,g7490,g2555);
	nand 	XG3498 	(g12147,g8201,g8302);
	nand 	XG3499 	(g11993,g8302,g1894);
	nand 	XG3500 	(g12188,g1894,g8249);
	nor 	XG3501 	(g12432,g8249,g1894);
	or 	XG3502 	(g8790,I12783,I12782);
	and 	XG3503 	(I24030,g3396,g8016,g8390);
	and 	XG3504 	(I24018,g3396,g8390,g8155);
	nor 	XG3505 	(g11357,g8561,g8558);
	not 	XG3506 	(g11043,g8561);
	not 	XG3507 	(g10357,g6825);
	nand 	XG3508 	(g10726,g1061,g979,g7661,g7304);
	nand 	XG3509 	(I12076,I12074,g979);
	not 	XG3510 	(g10368,g6887);
	nand 	XG3511 	(I14257,g3133,g8154);
	nand 	XG3512 	(g12413,g5654,g7521);
	nand 	XG3513 	(I13183,I13182,g6500);
	nand 	XG3514 	(I11865,I11864,g4434);
	nor 	XG3515 	(g12198,g9800,g9797);
	and 	XG3516 	(g11035,g9800,g5441);
	and 	XG3517 	(I24524,g9716,g5046,g5041);
	and 	XG3518 	(I13937,g7261,g7293,g7340);
	not 	XG3519 	(g10395,g6995);
	nand 	XG3520 	(I13565,I13564,g2648);
	nand 	XG3521 	(g12151,g8211,g8316);
	nand 	XG3522 	(g11975,g8316,g8267);
	nand 	XG3523 	(g12119,g8267,g2351);
	nand 	XG3524 	(g11117,g8239,g8186,g8087);
	not 	XG3525 	(g9772,I13352);
	nand 	XG3526 	(g12014,g703,g7197);
	nand 	XG3527 	(g12042,g703,g9086);
	nor 	XG3528 	(g11309,g8728,g8587);
	not 	XG3529 	(g11753,g8587);
	not 	XG3530 	(g8542,I12644);
	and 	XG3531 	(g10724,g8728,g3689);
	nand 	XG3532 	(I13731,I13729,g4537);
	not 	XG3533 	(g7626,I12112);
	nand 	XG3534 	(I13750,I13749,g4608);
	nor 	XG3535 	(g10555,g4608,g4601,g7227);
	not 	XG3536 	(g10374,g6903);
	not 	XG3537 	(g11741,g10033);
	nand 	XG3538 	(I14480,g655,g10074);
	nand 	XG3539 	(g12197,g5290,g7296);
	not 	XG3540 	(g10107,I13606);
	nand 	XG3541 	(I13079,I13077,g5467);
	not 	XG3542 	(g6868,I11688);
	and 	XG3543 	(I14225,g262,g8406,g255,g8457);
	nand 	XG3544 	(I13443,I13442,g262);
	nor 	XG3545 	(g12017,g9586,g9969);
	nand 	XG3546 	(g11445,g3976,g9771);
	nand 	XG3547 	(I13463,I13462,g2380);
	nor 	XG3548 	(g12246,g9883,g9880);
	not 	XG3549 	(g11866,g9883);
	nor 	XG3550 	(g10831,g7827,g7690);
	nand 	XG3551 	(g11396,g4688,g8713);
	nand 	XG3552 	(g12196,g4688,g8764);
	not 	XG3553 	(g10351,g6802);
	nand 	XG3554 	(g12227,g8330,g8418);
	nand 	XG3555 	(g12053,g8418,g2587);
	nand 	XG3556 	(g12287,g2587,g8381);
	nor 	XG3557 	(g12540,g8381,g2587);
	not 	XG3558 	(g8135,I12418);
	not 	XG3559 	(I14046,g9900);
	and 	XG3560 	(I24003,g3045,g8334,g8097);
	and 	XG3561 	(I24015,g3045,g7975,g8334);
	nand 	XG3562 	(g12341,g5308,g7512);
	not 	XG3563 	(g6976,I11750);
	not 	XG3564 	(g11030,g8292);
	not 	XG3565 	(g10389,g6986);
	not 	XG3566 	(g10386,g6982);
	nand 	XG3567 	(I12075,I12074,g996);
	and 	XG3568 	(g11028,g5428,g9730);
	nand 	XG3569 	(g12317,g6486,g10026);
	nand 	XG3570 	(I12469,I12468,g405);
	or 	XG3571 	(g8417,I12583,g1116,g1056);
	nand 	XG3572 	(g10909,g1116,g7304);
	nand 	XG3573 	(g10905,g7304,g1116);
	nor 	XG3574 	(g12204,g10160,g9927);
	not 	XG3575 	(g12804,g9927);
	not 	XG3576 	(g9864,I13424);
	and 	XG3577 	(g11114,g10160,g5689);
	nor 	XG3578 	(g12443,g9300,g9374);
	not 	XG3579 	(g12738,g9374);
	nor 	XG3580 	(g12772,g9300,g5188);
	nand 	XG3581 	(I12279,I12277,g1472);
	and 	XG3582 	(g12812,g9158,g518);
	nand 	XG3583 	(I14185,g3470,g8442);
	nor 	XG3584 	(g11584,g8172,g8229);
	not 	XG3585 	(g11754,g8229);
	nor 	XG3586 	(g11763,g8172,g3881);
	nor 	XG3587 	(g12467,g9407,g9472);
	nor 	XG3588 	(g12806,g9407,g9472);
	nor 	XG3589 	(g12755,g9407,g6555);
	nand 	XG3590 	(g10951,g7868,g7845);
	not 	XG3591 	(I15250,g9152);
	not 	XG3592 	(g12779,g9444);
	nand 	XG3593 	(I15087,g2393,g9832);
	nor 	XG3594 	(g10695,g8407,g8462);
	nor 	XG3595 	(g10649,g8407,g1183);
	nand 	XG3596 	(g12024,g8418,g8381);
	nand 	XG3597 	(g12195,g8381,g2619);
	not 	XG3598 	(g12122,g9705);
	not 	XG3599 	(g7632,I12117);
	nor 	XG3600 	(g11885,g7167,g7153);
	not 	XG3601 	(g10402,g7023);
	not 	XG3602 	(g12018,g9538);
	nand 	XG3603 	(g11245,g7697,g7733,g7636);
	not 	XG3604 	(I13979,g7733);
	not 	XG3605 	(g8778,I12758);
	not 	XG3606 	(g6971,I11737);
	not 	XG3607 	(g6789,I11635);
	not 	XG3608 	(I14550,g10072);
	nand 	XG3609 	(I12402,I12401,g3808);
	nand 	XG3610 	(I13383,I13382,g269);
	not 	XG3611 	(g10376,g6923);
	not 	XG3612 	(g12295,g7139);
	nor 	XG3613 	(g11276,g8691,g8534);
	not 	XG3614 	(g11735,g8534);
	not 	XG3615 	(g8481,I12618);
	and 	XG3616 	(g10706,g8691,g3338);
	not 	XG3617 	(g10371,g6918);
	not 	XG3618 	(g10373,g6917);
	not 	XG3619 	(g11042,g8691);
	nor 	XG3620 	(g11563,g8011,g8059);
	nor 	XG3621 	(g11473,g8059,g8107);
	nor 	XG3622 	(g11435,g3171,g8107);
	nor 	XG3623 	(g12571,g9451,g9511);
	not 	XG3624 	(g12805,g9511);
	nor 	XG3625 	(g12824,g9451,g5881);
	nand 	XG3626 	(g11446,g8734,g6941,g8700);
	not 	XG3627 	(g10375,g6941);
	and 	XG3628 	(g10898,g9100,g3706);
	nand 	XG3629 	(g12185,g799,g9905);
	not 	XG3630 	(g7993,I12333);
	not 	XG3631 	(g6767,I11626);
	not 	XG3632 	(I14455,g10197);
	not 	XG3633 	(g11812,g7567);
	not 	XG3634 	(g10881,g7567);
	not 	XG3635 	(g10872,g7567);
	not 	XG3636 	(g10621,g7567);
	nand 	XG3637 	(I13066,I13065,g4308);
	and 	XG3638 	(g10674,g2130,g10200,g6841);
	and 	XG3639 	(g10719,g2130,g2138,g6841);
	not 	XG3640 	(g7623,I12103);
	nand 	XG3641 	(g10610,g7490,g7462);
	and 	XG3642 	(g11978,g7462,g2629);
	and 	XG3643 	(I24546,g9716,g5052,g5046);
	nand 	XG3644 	(g10566,g7356,g7315);
	nand 	XG3645 	(g11992,g1772,g7275);
	nand 	XG3646 	(g10618,g9913,g10153);
	not 	XG3647 	(g10370,g7095);
	nand 	XG3648 	(I13499,I13497,g232);
	not 	XG3649 	(g10411,g7086);
	nand 	XG3650 	(g11190,g3447,g8539);
	not 	XG3651 	(g6973,I11743);
	nand 	XG3652 	(I11879,I11877,g4430);
	not 	XG3653 	(I15205,g10139);
	not 	XG3654 	(g10273,I13708);
	nand 	XG3655 	(I11878,I11877,g4388);
	not 	XG3656 	(g8470,I12605);
	not 	XG3657 	(I14409,g8364);
	not 	XG3658 	(g8572,I12654);
	nor 	XG3659 	(g11119,g9203,g9180);
	not 	XG3660 	(g8032,I12355);
	not 	XG3661 	(g7121,I11820);
	nor 	XG3662 	(g11666,g8125,g8172);
	not 	XG3663 	(g11884,g8125);
	nand 	XG3664 	(I13110,I13109,g5808);
	not 	XG3665 	(g10406,g7046);
	nand 	XG3666 	(g12125,g5101,g9728);
	nor 	XG3667 	(g12081,g9694,g10079);
	or 	XG3668 	(g10800,g952,g7517);
	nand 	XG3669 	(g11200,g3798,g8592);
	not 	XG3670 	(g10397,g7018);
	not 	XG3671 	(I15223,g10119);
	nand 	XG3672 	(I15002,g1700,g9691);
	not 	XG3673 	(g10361,g6841);
	not 	XG3674 	(g10366,g6895);
	nand 	XG3675 	(I13519,I13518,g2514);
	not 	XG3676 	(g8795,I12793);
	not 	XG3677 	(g10396,g6997);
	nor 	XG3678 	(g12046,g9640,g10036);
	not 	XG3679 	(I14119,g7824);
	not 	XG3680 	(g10405,g7064);
	not 	XG3681 	(I14593,g9978);
	not 	XG3682 	(g6856,I11682);
	and 	XG3683 	(g11427,g7158,g5706);
	nand 	XG3684 	(g11544,g4045,g3990,g8700);
	not 	XG3685 	(g8405,I12572);
	or 	XG3686 	(g8921,I12903,I12902);
	nand 	XG3687 	(I12841,I12840,g4222);
	not 	XG3688 	(g7148,I11835);
	nor 	XG3689 	(g11231,g4793,g4801,g7928);
	nor 	XG3690 	(g11261,g9030,g4801,g7928);
	not 	XG3691 	(I13968,g7697);
	not 	XG3692 	(g8757,I12746);
	not 	XG3693 	(g10541,g9407);
	nand 	XG3694 	(g11134,g8301,g8240,g8138);
	not 	XG3695 	(g10897,g7601);
	not 	XG3696 	(g11849,g7601);
	not 	XG3697 	(g10652,g7601);
	not 	XG3698 	(g10882,g7601);
	not 	XG3699 	(g12823,g9206);
	not 	XG3700 	(g11413,g9100);
	nand 	XG3701 	(I12263,I12261,g1448);
	nor 	XG3702 	(g11907,g7184,g7170);
	not 	XG3703 	(I14862,g8092);
	not 	XG3704 	(g6832,I11665);
	not 	XG3705 	(g7766,I12189);
	nor 	XG3706 	(g12659,g9392,g9451);
	not 	XG3707 	(g10540,g9392);
	nor 	XG3708 	(g11976,g7379,g9595);
	not 	XG3709 	(g12051,g9595);
	nand 	XG3710 	(g12192,g2319,g8267);
	nor 	XG3711 	(g12437,g8267,g2319);
	not 	XG3712 	(g9687,I13287);
	nand 	XG3713 	(g12255,g6140,g9958);
	and 	XG3714 	(g10966,g7948,g9226);
	nand 	XG3715 	(g11149,g7948,g1564);
	not 	XG3716 	(g10980,g9051);
	not 	XG3717 	(g11513,g7948);
	not 	XG3718 	(g11786,g7549);
	not 	XG3719 	(g12233,g10338);
	nand 	XG3720 	(g12008,g5798,g9932);
	nand 	XG3721 	(I13751,I13749,g4584);
	not 	XG3722 	(g10142,I13637);
	not 	XG3723 	(I14537,g10106);
	not 	XG3724 	(g6782,I11632);
	not 	XG3725 	(g11841,g9800);
	not 	XG3726 	(g8038,I12360);
	not 	XG3727 	(g8812,I12805);
	not 	XG3728 	(I13990,g7636);
	not 	XG3729 	(g10392,g6989);
	not 	XG3730 	(g8763,I12749);
	not 	XG3731 	(g10381,g6957);
	not 	XG3732 	(g11889,g9954);
	not 	XG3733 	(I14823,g8056);
	not 	XG3734 	(g6821,I11655);
	not 	XG3735 	(g8411,I12577);
	not 	XG3736 	(g7633,I12120);
	or 	XG3737 	(g12768,g7202,g7785);
	not 	XG3738 	(g10795,g7202);
	not 	XG3739 	(g12345,g7158);
	not 	XG3740 	(g7634,I12123);
	or 	XG3741 	(g8476,I12611,g1459,g1399);
	nand 	XG3742 	(g12307,g5983,g7395);
	nand 	XG3743 	(I12850,I12848,g4277);
	nand 	XG3744 	(I12849,I12848,g4281);
	not 	XG3745 	(g11815,g7582);
	nand 	XG3746 	(g12428,g6358,g7472);
	not 	XG3747 	(g10393,g6991);
	not 	XG3748 	(g7196,I11860);
	nand 	XG3749 	(I13141,I13139,g6159);
	not 	XG3750 	(g10960,g9007);
	and 	XG3751 	(g10917,g1087,g9174);
	not 	XG3752 	(g10518,g9311);
	not 	XG3753 	(g7738,I12176);
	and 	XG3754 	(g12135,g9959,g9684);
	not 	XG3755 	(g6928,I11716);
	not 	XG3756 	(g6888,I11701);
	nand 	XG3757 	(g11892,g9086,g7777);
	nor 	XG3758 	(g11999,g7423,g9654);
	nand 	XG3759 	(g10551,g7356,g1728);
	not 	XG3760 	(g11714,g8107);
	not 	XG3761 	(g12054,g7690);
	not 	XG3762 	(g10708,g7836);
	not 	XG3763 	(g10414,g7092);
	not 	XG3764 	(g8357,I12538);
	nor 	XG3765 	(g11039,g9092,g9056);
	and 	XG3766 	(g11083,g802,g8836);
	nand 	XG3767 	(g11679,g802,g8836);
	nand 	XG3768 	(g12464,g10191,g7087,g10169);
	and 	XG3769 	(g11496,g7495,g4382);
	not 	XG3770 	(g10407,g7063);
	not 	XG3771 	(g11811,g9724);
	not 	XG3772 	(g10323,I13744);
	not 	XG3773 	(g11861,g8070);
	not 	XG3774 	(g10420,g9239);
	not 	XG3775 	(g9155,I12997);
	nand 	XG3776 	(I13730,I13729,g4534);
	not 	XG3777 	(g8740,I12735);
	nor 	XG3778 	(g11493,g8967,g8964);
	and 	XG3779 	(g10856,g8967,g4269);
	not 	XG3780 	(g11031,g8609);
	not 	XG3781 	(g10359,g6830);
	not 	XG3782 	(g6955,I11726);
	nor 	XG3783 	(g10893,g7749,g7715,g1189);
	not 	XG3784 	(g10390,g6987);
	not 	XG3785 	(g7994,I12336);
	not 	XG3786 	(g11344,g9015);
	and 	XG3787 	(g12284,g7557,g1532);
	nor 	XG3788 	(g10918,g7778,g7751,g1532);
	not 	XG3789 	(g11736,g8165);
	not 	XG3790 	(g10497,g10102);
	not 	XG3791 	(g10061,I13581);
	not 	XG3792 	(g10369,g6873);
	not 	XG3793 	(g10400,g7002);
	nand 	XG3794 	(g10961,g7876,g1442);
	nor 	XG3795 	(g11363,g8751,g8626);
	not 	XG3796 	(g11122,g8751);
	not 	XG3797 	(g10372,g6900);
	not 	XG3798 	(g7617,I12089);
	nand 	XG3799 	(g11971,g8302,g8249);
	nand 	XG3800 	(g11955,g1917,g8302);
	nor 	XG3801 	(g12189,g8302,g1917);
	nand 	XG3802 	(I12218,I12217,g1437);
	nand 	XG3803 	(g12073,g6490,g10058);
	nand 	XG3804 	(g11251,g3092,g8438);
	nor 	XG3805 	(g12166,g10124,g9856);
	not 	XG3806 	(g11865,g10124);
	not 	XG3807 	(g7526,I12013);
	not 	XG3808 	(g7502,I11992);
	not 	XG3809 	(g8134,I12415);
	not 	XG3810 	(g12086,g9654);
	not 	XG3811 	(g10378,g6926);
	not 	XG3812 	(g10353,g6803);
	not 	XG3813 	(g7660,I12144);
	not 	XG3814 	(g12778,g9856);
	not 	XG3815 	(g9780,I13360);
	not 	XG3816 	(g7074,I11801);
	not 	XG3817 	(g10410,g7069);
	nand 	XG3818 	(I12205,I12203,g1135);
	not 	XG3819 	(g11721,g10074);
	not 	XG3820 	(g10216,I13684);
	not 	XG3821 	(g10399,g7017);
	not 	XG3822 	(g6977,I11753);
	not 	XG3823 	(g6867,I11685);
	not 	XG3824 	(g10230,I13694);
	nand 	XG3825 	(I12346,I12344,g3111);
	not 	XG3826 	(g11927,g10207);
	nor 	XG3827 	(g11385,g7985,g8021);
	nor 	XG3828 	(g11692,g7985,g8021);
	not 	XG3829 	(g11796,g7985);
	nor 	XG3830 	(g11658,g3506,g8021);
	not 	XG3831 	(g7616,I12086);
	not 	XG3832 	(g10409,g7087);
	nand 	XG3833 	(g12245,g5637,g7344);
	not 	XG3834 	(I14570,g7932);
	not 	XG3835 	(g12440,g9985);
	not 	XG3836 	(g8971,I12927);
	nand 	XG3837 	(g12369,g637,g9049);
	not 	XG3838 	(g11214,g9602);
	not 	XG3839 	(g11779,g9602);
	not 	XG3840 	(g7791,I12199);
	nor 	XG3841 	(g12708,g9462,g9518);
	not 	XG3842 	(g10564,g9462);
	not 	XG3843 	(g12047,g9591);
	not 	XG3844 	(g10725,g7846);
	not 	XG3845 	(g11810,g9664);
	not 	XG3846 	(g11233,g9664);
	not 	XG3847 	(g10350,g6800);
	not 	XG3848 	(g11472,g7918);
	not 	XG3849 	(g7689,I12159);
	not 	XG3850 	(g7593,I12061);
	not 	XG3851 	(g11110,g8728);
	not 	XG3852 	(g10404,g7026);
	not 	XG3853 	(g10394,g6994);
	nand 	XG3854 	(I13510,I13509,g2089);
	not 	XG3855 	(g10408,g7049);
	not 	XG3856 	(g7516,I12003);
	not 	XG3857 	(g11316,g8967);
	nand 	XG3858 	(I12097,I12096,g1339);
	not 	XG3859 	(g10412,g7072);
	nand 	XG3860 	(I11825,I11824,g4593);
	not 	XG3861 	(g11038,g8632);
	nand 	XG3862 	(I12373,I12372,g3457);
	not 	XG3863 	(g10295,I13723);
	not 	XG3864 	(g11832,g8011);
	not 	XG3865 	(g7527,I12016);
	not 	XG3866 	(g10352,g6804);
	not 	XG3867 	(g11888,g10160);
	not 	XG3868 	(g11762,g7964);
	not 	XG3869 	(g11910,g10185);
	not 	XG3870 	(g7625,I12109);
	not 	XG3871 	(g10382,g6958);
	not 	XG3872 	(g8880,I12861);
	not 	XG3873 	(g11011,g10274);
	not 	XG3874 	(g7648,I12135);
	and 	XG3875 	(g12259,g640,g9480);
	nand 	XG3876 	(g12323,g640,g9480);
	not 	XG3877 	(g8595,I12666);
	not 	XG3878 	(g11769,g8626);
	and 	XG3879 	(I24505,g5057,g9229,g9607);
	and 	XG3880 	(I24482,g5057,g9607,g9364);
	and 	XG3881 	(g10736,g8751,g4040);
	nand 	XG3882 	(I13111,I13109,g5813);
	and 	XG3883 	(g11915,g7315,g1802);
	nor 	XG3884 	(g12581,g6219,g9569);
	nand 	XG3885 	(g12111,g9166,g847);
	nand 	XG3886 	(g11951,g703,g847,g9166);
	nor 	XG3887 	(g11621,g7985,g3512);
	nand 	XG3888 	(I12842,I12840,g4235);
	nand 	XG3889 	(I15212,g1714,g10035);
	nand 	XG3890 	(g11443,g3649,g9916);
	nand 	XG3891 	(g11411,g3625,g9713);
	nor 	XG3892 	(g11610,g3155,g7980);
	and 	XG3893 	(g10883,g9061,g3355);
	nand 	XG3894 	(I15078,g1968,g9827);
	nand 	XG3895 	(g10511,g4621,g7202,g4628);
	nand 	XG3896 	(g11320,g7202,g4621,g4633);
	and 	XG3897 	(g11967,g7802,g311);
	nor 	XG3898 	(g11252,g3057,g8620);
	nor 	XG3899 	(g11191,g9030,g4801,g4776);
	nor 	XG3900 	(g11213,g9030,g7892,g4776);
	nand 	XG3901 	(g11155,g9030,g7892,g4776);
	nor 	XG3902 	(g10510,g4584,g4593,g7183);
	nor 	XG3903 	(g10803,g7503,g1384);
	nor 	XG3904 	(g10821,g1384,g7503);
	nor 	XG3905 	(g12405,g5180,g9374);
	and 	XG3906 	(g10822,g8514,g4264);
	nand 	XG3907 	(g11489,g3618,g9661);
	nand 	XG3908 	(g12207,g5794,g9887);
	nand 	XG3909 	(g12035,g6144,g10000);
	nand 	XG3910 	(I12403,I12401,g3813);
	and 	XG3911 	(g10896,g8654,g1205);
	and 	XG3912 	(I24616,g9946,g6088,g6082);
	nand 	XG3913 	(g10929,g7854,g1099);
	nand 	XG3914 	(g12232,g4878,g8804);
	nand 	XG3915 	(g11426,g4878,g8742);
	nand 	XG3916 	(g12343,g5630,g7470);
	nand 	XG3917 	(g12459,g5623,g7437);
	nand 	XG3918 	(g12115,g8249,g1926);
	nand 	XG3919 	(g11674,g4674,g8676);
	nand 	XG3920 	(g12124,g4674,g8741);
	nand 	XG3921 	(g12521,g5969,g7471);
	nand 	XG3922 	(g12356,g6012,g7438);
	nand 	XG3923 	(g10567,g7405,g1862);
	nor 	XG3924 	(g11932,g9166,g843);
	nand 	XG3925 	(g12306,g5666,g7394);
	nand 	XG3926 	(g12588,g6386,g6336,g10169);
	nand 	XG3927 	(g12463,g6322,g7513);
	nand 	XG3928 	(g12587,g6315,g7497);
	nand 	XG3929 	(g12159,g4864,g8765);
	nand 	XG3930 	(g11707,g4864,g8718);
	and 	XG3931 	(g12186,g7519,g1178);
	and 	XG3932 	(g10878,g1135,g7858);
	and 	XG3933 	(I24051,g8492,g3385,g3380);
	and 	XG3934 	(g11044,g10124,g5343);
	nand 	XG3935 	(g11312,g3794,g8565);
	nand 	XG3936 	(g12152,g8324,g2485);
	and 	XG3937 	(g10829,g4375,g7289);
	and 	XG3938 	(g11546,g4375,g7289);
	nand 	XG3939 	(g11639,g4722,g8933);
	nand 	XG3940 	(g12589,g6692,g7591);
	nand 	XG3941 	(g12525,g6668,g7522);
	nand 	XG3942 	(I13140,I13139,g6154);
	and 	XG3943 	(g10528,g9051,g1576);
	nand 	XG3944 	(g12080,g8201,g1917);
	and 	XG3945 	(I24048,g8426,g3040,g3034);
	nand 	XG3946 	(g11543,g3969,g9714);
	nand 	XG3947 	(g11424,g4012,g9662);
	and 	XG3948 	(g10501,g9007,g1233);
	nand 	XG3949 	(g12357,g6329,g7439);
	nor 	XG3950 	(g12288,g8418,g2610);
	nand 	XG3951 	(g12153,g8330,g2610);
	nand 	XG3952 	(g12000,g2610,g8418);
	and 	XG3953 	(g11397,g7139,g5360);
	nand 	XG3954 	(I12262,I12261,g1454);
	or 	XG3955 	(g10802,g1296,g7533);
	and 	XG3956 	(g11163,g10224,g6727);
	nor 	XG3957 	(g11747,g8114,g3530);
	nand 	XG3958 	(I13067,I13065,g4304);
	nand 	XG3959 	(g11858,g3010,g9014);
	and 	XG3960 	(g12219,g7532,g1189);
	nand 	XG3961 	(g10569,g7418,g2287);
	nor 	XG3962 	(g10793,g7503,g1389);
	nand 	XG3963 	(I14923,g5835,g9558);
	nor 	XG3964 	(g10666,g1171,g8462);
	nor 	XG3965 	(g11248,g4983,g4991,g7953);
	nand 	XG3966 	(g11394,g3661,g9600);
	nand 	XG3967 	(g11442,g3343,g3288,g8644);
	and 	XG3968 	(g11497,g7192,g6398);
	nand 	XG3969 	(I15051,g2259,g9759);
	nand 	XG3970 	(g10928,g417,g8137,g8181);
	nor 	XG3971 	(g10709,g351,g7499);
	nor 	XG3972 	(g12651,g5511,g9269);
	and 	XG3973 	(g11019,g9036,g5092);
	and 	XG3974 	(I24579,g9875,g5736,g5731);
	and 	XG3975 	(I24597,g9875,g5742,g5736);
	nand 	XG3976 	(g12052,g2465,g7387);
	nand 	XG3977 	(g11326,g370,g365,g376,g8993);
	nor 	XG3978 	(g11729,g8059,g3179);
	nand 	XG3979 	(I14289,g3835,g8282);
	and 	XG3980 	(g12761,g7567,g969);
	and 	XG3981 	(g10616,g174,g7998);
	nand 	XG3982 	(I12242,I12240,g1105);
	and 	XG3983 	(g10890,g1105,g7858);
	nor 	XG3984 	(g12193,g8316,g2342);
	nand 	XG3985 	(g11959,g2342,g8316);
	nand 	XG3986 	(g12084,g8211,g2342);
	nand 	XG3987 	(g11395,g3983,g9601);
	nand 	XG3988 	(g12340,g8984,g4888);
	and 	XG3989 	(g11016,g8984,g4888);
	nand 	XG3990 	(g10935,g7352,g1459);
	nand 	XG3991 	(g10939,g1459,g7352);
	nand 	XG3992 	(g10561,g5712,g7157);
	and 	XG3993 	(I24067,g8553,g3736,g3731);
	and 	XG3994 	(I24075,g8553,g3742,g3736);
	and 	XG3995 	(g11037,g9184,g6128);
	nand 	XG3996 	(I13384,I13382,g246);
	and 	XG3997 	(g11024,g9070,g5436);
	nand 	XG3998 	(I13444,I13442,g239);
	nand 	XG3999 	(g10515,g5022,g10337);
	nand 	XG4000 	(g11491,g4000,g9982);
	and 	XG4001 	(g10947,g1430,g9200);
	and 	XG4002 	(I14198,g8180,g232,g8237,g225);
	nor 	XG4003 	(g12515,g5873,g9511);
	nand 	XG4004 	(g11997,g8316,g2319);
	nand 	XG4005 	(I14788,g6167,g9891);
	nand 	XG4006 	(g12087,g2599,g7431);
	and 	XG4007 	(g10967,g1448,g7880);
	nand 	XG4008 	(g11903,g3712,g9099);
	nor 	XG4009 	(g12593,g5164,g9234);
	nor 	XG4010 	(g12785,g6549,g9472);
	nand 	XG4011 	(I12278,I12277,g1467);
	nand 	XG4012 	(g12522,g6040,g5990,g10133);
	and 	XG4013 	(g10675,g8500,g3436);
	and 	XG4014 	(g11045,g9883,g5787);
	and 	XG4015 	(g10704,g2130,g10200,g2145);
	nor 	XG4016 	(g11184,g9040,g513);
	nand 	XG4017 	(g12412,g5348,g5297,g10044);
	nor 	XG4018 	(g12208,g5759,g10096);
	nor 	XG4019 	(g11537,g3873,g8229);
	nand 	XG4020 	(g11356,g3632,g9552);
	nor 	XG4021 	(g10801,g7479,g1041);
	nor 	XG4022 	(g10819,g1041,g7479);
	nand 	XG4023 	(g11979,g5452,g9861);
	nor 	XG4024 	(g11306,g8647,g3412);
	and 	XG4025 	(I24549,g9792,g5390,g5385);
	and 	XG4026 	(I24027,g8426,g3034,g3029);
	and 	XG4027 	(g10707,g8561,g3787);
	nor 	XG4028 	(g11891,g9166,g812);
	nand 	XG4029 	(g11302,g3281,g9496);
	nand 	XG4030 	(g11490,g3694,g3639,g8666);
	nand 	XG4031 	(g11961,g5105,g9777);
	nor 	XG4032 	(g11313,g3759,g8669);
	nor 	XG4033 	(g12371,g8195,g1760);
	nand 	XG4034 	(g11970,g8241,g1760);
	nand 	XG4035 	(g12145,g1760,g8195);
	nand 	XG4036 	(g12293,g5283,g7436);
	nand 	XG4037 	(g12411,g5276,g7393);
	nand 	XG4038 	(I13566,I13564,g2652);
	nand 	XG4039 	(I14516,g661,g10147);
	nor 	XG4040 	(g12798,g9381,g5535);
	nand 	XG4041 	(g10916,g7854,g1146);
	and 	XG4042 	(I24064,g8492,g3391,g3385);
	and 	XG4043 	(g10999,g1472,g7880);
	and 	XG4044 	(g11937,g7362,g1936);
	nor 	XG4045 	(g12591,g9040,g504);
	nand 	XG4046 	(g12169,g5448,g9804);
	and 	XG4047 	(g11036,g5774,g9806);
	and 	XG4048 	(I24576,g9792,g5396,g5390);
	and 	XG4049 	(g11893,g7268,g1668);
	nor 	XG4050 	(g12711,g9326,g6209);
	nand 	XG4051 	(g11990,g703,g9166);
	and 	XG4052 	(g11740,g703,g8769);
	nand 	XG4053 	(g10583,g862,g7475);
	nand 	XG4054 	(g11002,g862,g7475);
	nand 	XG4055 	(I13850,g7397,g862);
	nand 	XG4056 	(g12048,g2040,g7369);
	nand 	XG4057 	(I14228,g8055,g979);
	and 	XG4058 	(g10676,g3774,g8506);
	and 	XG4059 	(I24600,g9946,g6082,g6077);
	nor 	XG4060 	(g10671,g8466,g1526);
	nor 	XG4061 	(g12662,g9274,g5863);
	nand 	XG4062 	(g11675,g4912,g8984);
	nand 	XG4063 	(g10552,g7374,g2153);
	or 	XG4064 	(g11370,g550,g8807);
	and 	XG4065 	(g10948,g1478,g7880);
	and 	XG4066 	(g10619,g7907,g3080);
	nor 	XG4067 	(g11669,g8026,g3863);
	nand 	XG4068 	(I13454,I13452,g1959);
	nand 	XG4069 	(g12120,g8273,g2476);
	nor 	XG4070 	(g12729,g8139,g1657);
	nand 	XG4071 	(g12044,g8139,g1657);
	nand 	XG4072 	(g11676,g385,g376,g8944,g358);
	and 	XG4073 	(g10655,g3423,g8440);
	nand 	XG4074 	(g12429,g6675,g7473);
	nand 	XG4075 	(I12546,I12544,g194);
	nor 	XG4076 	(g11755,g8796,g4709);
	nand 	XG4077 	(g11409,g3298,g9842);
	and 	XG4078 	(g12527,g667,g8680);
	nand 	XG4079 	(I14733,g5475,g9732);
	nand 	XG4080 	(g12639,g6732,g6682,g10194);
	nand 	XG4081 	(I15121,g2102,g9910);
	nor 	XG4082 	(g12150,g8259,g2208);
	nand 	XG4083 	(g12049,g8150,g2208);
	nand 	XG4084 	(g11938,g2208,g8259);
	nor 	XG4085 	(g10899,g8451,g4064);
	and 	XG4086 	(g10657,g4064,g8451);
	nor 	XG4087 	(g11780,g8822,g4899);
	nand 	XG4088 	(I13045,I13043,g5120);
	nand 	XG4089 	(I15363,g2675,g10182);
	and 	XG4090 	(I24619,g10014,g6428,g6423);
	and 	XG4091 	(I24625,g10014,g6434,g6428);
	and 	XG4092 	(g11116,g6466,g9960);
	nand 	XG4093 	(I13392,I13390,g1825);
	nand 	XG4094 	(g11974,g8259,g2185);
	nand 	XG4095 	(I15306,g2407,g10116);
	nor 	XG4096 	(g12146,g8241,g1783);
	nand 	XG4097 	(g11936,g1783,g8241);
	and 	XG4098 	(g10902,g1129,g7858);
	and 	XG4099 	(g11916,g7328,g2227);
	nand 	XG4100 	(I13402,I13401,g2246);
	nor 	XG4101 	(g12333,g8139,g1624);
	nand 	XG4102 	(g12112,g1624,g8139);
	and 	XG4103 	(g10720,g2689,g10219,g2704);
	and 	XG4104 	(g10732,g2689,g2697,g6850);
	and 	XG4105 	(g10705,g2689,g10219,g6850);
	nor 	XG4106 	(g10491,g9576,g6573);
	nor 	XG4107 	(g12479,g8310,g2028);
	nand 	XG4108 	(g12020,g8365,g2028);
	nand 	XG4109 	(g12222,g2028,g8310);
	and 	XG4110 	(g10925,g956,g7858);
	nand 	XG4111 	(g11381,g3274,g9660);
	nand 	XG4112 	(g12460,g5694,g5644,g10093);
	and 	XG4113 	(g12730,g4349,g9024);
	nand 	XG4114 	(I15298,g1982,g10112);
	nand 	XG4115 	(g12638,g6661,g7514);
	nand 	XG4116 	(I14853,g5142,g9433);
	nor 	XG4117 	(g12223,g8365,g2051);
	nand 	XG4118 	(g11973,g2051,g8365);
	nor 	XG4119 	(g11280,g3408,g8647);
	nand 	XG4120 	(I13335,I13334,g1687);
	nand 	XG4121 	(I14169,g3119,g8389);
	nor 	XG4122 	(g12847,g10430,g6838);
	nor 	XG4123 	(g12850,g6845,g10430);
	nor 	XG4124 	(g12848,g10430,g6839);
	nor 	XG4125 	(g12855,g6854,g10430);
	nor 	XG4126 	(g12856,g6855,g10430);
	nor 	XG4127 	(g12852,g10430,g6847);
	nor 	XG4128 	(g12846,g10430,g6837);
	nor 	XG4129 	(g12854,g10430,g6849);
	nor 	XG4130 	(g12849,g10430,g6840);
	nor 	XG4131 	(g12853,g10430,g6848);
	nor 	XG4132 	(g12851,g10430,g6846);
	not 	XG4133 	(I15587,g11985);
	not 	XG4134 	(I15533,g11867);
	not 	XG4135 	(I15650,g12110);
	not 	XG4136 	(I15556,g11928);
	not 	XG4137 	(I15705,g12218);
	not 	XG4138 	(I15623,g12040);
	not 	XG4139 	(I15569,g11965);
	not 	XG4140 	(I15682,g12182);
	not 	XG4141 	(I15609,g12013);
	not 	XG4142 	(I15626,g12041);
	not 	XG4143 	(I15593,g11989);
	not 	XG4144 	(I16452,g11182);
	not 	XG4145 	(I15636,g12075);
	not 	XG4146 	(I16535,g11235);
	not 	XG4147 	(I15736,g12322);
	not 	XG4148 	(I15564,g11949);
	not 	XG4149 	(I16486,g11204);
	not 	XG4150 	(I15617,g12037);
	not 	XG4151 	(I15667,g12143);
	not 	XG4152 	(I16438,g11165);
	not 	XG4153 	(I15620,g12038);
	not 	XG4154 	(I15647,g12109);
	not 	XG4155 	(I15590,g11988);
	not 	XG4156 	(I15448,g10877);
	not 	XG4157 	(I15702,g12217);
	not 	XG4158 	(I15633,g12074);
	not 	XG4159 	(g13494,g11912);
	not 	XG4160 	(g13412,g11963);
	not 	XG4161 	(g13302,g12321);
	not 	XG4162 	(g13087,g12012);
	not 	XG4163 	(g13070,g11984);
	not 	XG4164 	(g13051,g11964);
	not 	XG4165 	(g14562,g12036);
	not 	XG4166 	(g14357,g12181);
	not 	XG4167 	(g14198,g12180);
	not 	XG4168 	(g14173,g12076);
	not 	XG4169 	(I15474,g10364);
	not 	XG4170 	(I16521,g10430);
	not 	XG4171 	(I15788,g10430);
	not 	XG4172 	(I16613,g10430);
	not 	XG4173 	(I16135,g10430);
	not 	XG4174 	(I15906,g10430);
	not 	XG4175 	(I15577,g10430);
	not 	XG4176 	(I16555,g10430);
	not 	XG4177 	(I16476,g10430);
	not 	XG4178 	(I15782,g10430);
	not 	XG4179 	(I15915,g10430);
	not 	XG4180 	(I15893,g10430);
	not 	XG4181 	(I16460,g10430);
	not 	XG4182 	(I16709,g10430);
	not 	XG4183 	(I16498,g10430);
	not 	XG4184 	(I16057,g10430);
	not 	XG4185 	(I16090,g10430);
	not 	XG4186 	(I15929,g10430);
	not 	XG4187 	(I16040,g10430);
	not 	XG4188 	(I15600,g10430);
	not 	XG4189 	(I16117,g10430);
	not 	XG4190 	(I16479,g10430);
	not 	XG4191 	(I15773,g10430);
	not 	XG4192 	(I16502,g10430);
	not 	XG4193 	(I15550,g10430);
	not 	XG4194 	(I16102,g10430);
	not 	XG4195 	(I16077,g10430);
	not 	XG4196 	(I16526,g10430);
	not 	XG4197 	(I16150,g10430);
	nor 	XG4198 	(g14415,g9590,g12147);
	and 	XG4199 	(g13081,g11122,g8626);
	not 	XG4200 	(g11631,g8595);
	nand 	XG4201 	(I15341,I15340,g10154);
	nand 	XG4202 	(g9391,I13111,I13110);
	nor 	XG4203 	(g14361,g9413,g12079);
	nand 	XG4204 	(g14940,g12581,g12744);
	nand 	XG4205 	(g14902,g12581,g7791);
	nand 	XG4206 	(g15036,g12581,g12780);
	nand 	XG4207 	(g12578,g10341,g7791);
	nand 	XG4208 	(g14861,g10341,g12744);
	nand 	XG4209 	(g15008,g10341,g12780);
	and 	XG4210 	(g10874,g6227,g6219,g7791);
	not 	XG4211 	(g11562,g7648);
	nor 	XG4212 	(g14178,g11083,g8899);
	nand 	XG4213 	(g14254,g11951,g11933,g11968);
	nor 	XG4214 	(g13336,g11011,g11330);
	not 	XG4215 	(g12885,g10382);
	nor 	XG4216 	(g11571,g3506,g3512,g10323);
	nand 	XG4217 	(g13955,g11527,g11621);
	nand 	XG4218 	(g13920,g11483,g11621);
	nor 	XG4219 	(g14094,g11083,g8770);
	not 	XG4220 	(g11470,g7625);
	nand 	XG4221 	(I14276,I14275,g8218);
	nand 	XG4222 	(I15193,g6005,g9935);
	and 	XG4223 	(I16671,g12415,g12461,g10185);
	nand 	XG4224 	(g8871,I12842,I12841);
	nor 	XG4225 	(g14313,g9250,g12016);
	and 	XG4226 	(g10733,g8542,g3625,g6905,g3639);
	nor 	XG4227 	(g11514,g3155,g3161,g10295);
	nand 	XG4228 	(g14008,g11435,g11610);
	nand 	XG4229 	(g14041,g11473,g11610);
	nand 	XG4230 	(g14234,g11881,g9177);
	nor 	XG4231 	(g13959,g11309,g3698);
	nand 	XG4232 	(g11533,g3698,g3639,g6905);
	nor 	XG4233 	(g14335,g9283,g12045);
	nand 	XG4234 	(I15147,g5659,g9864);
	or 	XG4235 	(g11372,g8038,g482,g490);
	not 	XG4236 	(g12835,g10352);
	nand 	XG4237 	(g14408,g11924,g6069);
	not 	XG4238 	(g11293,g7527);
	nor 	XG4239 	(g13913,g11083,g8859);
	nand 	XG4240 	(g14011,g11473,g10295);
	nand 	XG4241 	(g13980,g11435,g10295);
	nand 	XG4242 	(g8069,I12374,I12373);
	nand 	XG4243 	(g13291,g1500,g10715);
	or 	XG4244 	(g13006,g10034,g12284);
	or 	XG4245 	(g12982,g9968,g12220);
	nand 	XG4246 	(g13464,g4776,g4793,g10831);
	nand 	XG4247 	(g7133,I11826,I11825);
	not 	XG4248 	(g12909,g10412);
	nand 	XG4249 	(g7620,I12098,I12097);
	nand 	XG4250 	(g14758,g12405,g7704);
	nand 	XG4251 	(g14953,g12405,g12646);
	nand 	XG4252 	(g14656,g12405,g12553);
	nand 	XG4253 	(g14915,g10266,g12553);
	nand 	XG4254 	(g12402,g10266,g7704);
	nand 	XG4255 	(g14879,g10266,g12646);
	and 	XG4256 	(g10823,g5188,g5180,g7704);
	or 	XG4257 	(g13540,g10827,g10822);
	nor 	XG4258 	(g14124,g11083,g8830);
	not 	XG4259 	(g11269,g7516);
	not 	XG4260 	(g12905,g10408);
	nand 	XG4261 	(g9972,I13511,I13510);
	not 	XG4262 	(g12887,g10394);
	not 	XG4263 	(g12901,g10404);
	nand 	XG4264 	(g8124,I12403,I12402);
	not 	XG4265 	(g11401,g7593);
	not 	XG4266 	(g11677,g7689);
	or 	XG4267 	(g13662,g10917,g10896);
	nand 	XG4268 	(g13756,g12812,g203);
	nand 	XG4269 	(g13727,g12812,g168,g203,g174);
	nand 	XG4270 	(g13511,g12812,g203,g174,g182);
	nand 	XG4271 	(g13527,g12812,g203,g168,g182);
	not 	XG4272 	(g12839,g10350);
	nor 	XG4273 	(g13326,g10905,g10929);
	and 	XG4274 	(g14874,g10909,g1099);
	and 	XG4275 	(I16646,g12343,g12413,g10160);
	and 	XG4276 	(g11123,g9864,g5630,g7028,g5644);
	not 	XG4277 	(g12950,g12708);
	nand 	XG4278 	(g14943,g12622,g7791);
	nand 	XG4279 	(g14864,g10421,g7791);
	and 	XG4280 	(g14587,g10567,g10584);
	not 	XG4281 	(g10553,g8971);
	not 	XG4282 	(g11691,I14570);
	nor 	XG4283 	(g12101,g7074,g6336);
	nand 	XG4284 	(g12628,g6390,g6336,g7074);
	and 	XG4285 	(g11160,g10003,g6322,g7074,g6336);
	nor 	XG4286 	(g12173,g7074,g10050);
	not 	XG4287 	(g12902,g10409);
	not 	XG4288 	(g11429,g7616);
	nand 	XG4289 	(g14048,g11483,g11658);
	nand 	XG4290 	(g14075,g11527,g11658);
	nand 	XG4291 	(g14151,g11483,g11692);
	nand 	XG4292 	(g13923,g11527,g11692);
	not 	XG4293 	(g14192,g11385);
	nor 	XG4294 	(g14248,g10578,g6065);
	and 	XG4295 	(I16695,g12463,g12523,g10207);
	nand 	XG4296 	(g8010,I12346,I12345);
	not 	XG4297 	(I14964,g10230);
	not 	XG4298 	(g10365,g6867);
	not 	XG4299 	(g12891,g10399);
	not 	XG4300 	(I14939,g10216);
	nand 	XG4301 	(I14481,I14480,g10074);
	nand 	XG4302 	(g7803,I12205,I12204);
	not 	XG4303 	(g12904,g10410);
	and 	XG4304 	(g13541,g12308,g7069);
	not 	XG4305 	(g12749,g7074);
	not 	XG4306 	(g12497,g9780);
	not 	XG4307 	(I13857,g9780);
	and 	XG4308 	(g13492,g11865,g9856);
	not 	XG4309 	(g11609,g7660);
	nor 	XG4310 	(g14165,g11083,g8951);
	not 	XG4311 	(g12838,g10353);
	not 	XG4312 	(g12871,g10378);
	nand 	XG4313 	(I14713,I14712,g9671);
	not 	XG4314 	(g11181,g8134);
	and 	XG4315 	(g14097,g10632,g878);
	and 	XG4316 	(g14218,g10632,g875);
	nor 	XG4317 	(g13806,g4076,g11245);
	nor 	XG4318 	(g13831,g7666,g11245);
	nor 	XG4319 	(g14002,g11083,g8681);
	not 	XG4320 	(g11250,g7502);
	or 	XG4321 	(g13155,g11546,g11496);
	not 	XG4322 	(g11291,g7526);
	and 	XG4323 	(g11178,g10061,g6668,g7097,g6682);
	nand 	XG4324 	(g7823,I12219,I12218);
	nand 	XG4325 	(g9461,I13141,I13140);
	nand 	XG4326 	(I14249,I14247,g8091);
	and 	XG4327 	(g14612,g11993,g11971);
	not 	XG4328 	(g11430,g7617);
	nor 	XG4329 	(g13872,g11083,g8745);
	and 	XG4330 	(g14028,g11797,g8673);
	not 	XG4331 	(g12865,g10372);
	and 	XG4332 	(g13059,g11303,g6900);
	nand 	XG4333 	(g13288,g1442,g10946);
	nand 	XG4334 	(I15241,g6351,g10003);
	not 	XG4335 	(g12897,g10400);
	nand 	XG4336 	(g12941,g10537,g7167);
	nand 	XG4337 	(g7879,I12263,I12262);
	nand 	XG4338 	(g14177,g753,g11721,g11741);
	or 	XG4339 	(g14182,g753,g11721,g11741);
	not 	XG4340 	(g12866,g10369);
	or 	XG4341 	(g11025,g7831,g2980);
	not 	XG4342 	(g12721,g10061);
	and 	XG4343 	(g13567,g11948,g10102);
	nand 	XG4344 	(g13986,g11747,g10323);
	nand 	XG4345 	(g11480,g8906,g10323);
	and 	XG4346 	(g12692,g3530,g3522,g10323);
	not 	XG4347 	(g13322,g10918);
	nand 	XG4348 	(g9295,I13067,I13066);
	nor 	XG4349 	(g14417,g9648,g12149);
	nand 	XG4350 	(g13627,g8388,g11172);
	not 	XG4351 	(g11129,g7994);
	nand 	XG4352 	(g13834,g11773,g4754);
	and 	XG4353 	(g13345,g11773,g4754);
	not 	XG4354 	(g12883,g10390);
	not 	XG4355 	(g13314,g10893);
	and 	XG4356 	(g14589,g10569,g10586);
	and 	XG4357 	(g13265,g11493,g9018);
	not 	XG4358 	(g12843,g10359);
	nand 	XG4359 	(I15003,I15002,g9691);
	not 	XG4360 	(g13868,g11493);
	nand 	XG4361 	(I15088,I15087,g9832);
	nand 	XG4362 	(g13628,g11107,g3372);
	nand 	XG4363 	(g13486,g4966,g4983,g10862);
	nand 	XG4364 	(g13469,g10862,g4983);
	not 	XG4365 	(g12546,g8740);
	nor 	XG4366 	(g13954,g11276,g8663);
	nand 	XG4367 	(g10307,I13731,I13730);
	nand 	XG4368 	(g13000,g10598,g7228);
	and 	XG4369 	(g14061,g11834,g8715);
	not 	XG4370 	(g10608,g9155);
	nor 	XG4371 	(g12558,g5511,g5517,g7738);
	nand 	XG4372 	(g14848,g12453,g12651);
	nand 	XG4373 	(g14885,g12505,g12651);
	nand 	XG4374 	(g14051,g11527,g10323);
	nand 	XG4375 	(g14018,g11483,g10323);
	or 	XG4376 	(g13941,g11023,g11019);
	nand 	XG4377 	(g13909,g8803,g11674,g8847,g11396);
	nand 	XG4378 	(g14596,g9663,g12124,g9775,g12196);
	not 	XG4379 	(g12899,g10407);
	nor 	XG4380 	(g14867,g12314,g10191);
	not 	XG4381 	(g14232,g11083);
	not 	XG4382 	(g11236,g8357);
	nand 	XG4383 	(I15334,I15333,g10152);
	not 	XG4384 	(g12908,g10414);
	and 	XG4385 	(g13566,g12358,g7092);
	nand 	XG4386 	(I14510,I14508,g8721);
	nand 	XG4387 	(g14101,g11729,g11653);
	nand 	XG4388 	(g13873,g11729,g11566);
	nand 	XG4389 	(g14098,g8864,g11566);
	nand 	XG4390 	(g14069,g8864,g11653);
	and 	XG4391 	(g14566,g10551,g10566);
	nand 	XG4392 	(I14956,I14955,g9620);
	nand 	XG4393 	(g13911,g4917,g11834);
	and 	XG4394 	(g10828,g7640,g6888);
	not 	XG4395 	(g11702,g6928);
	nand 	XG4396 	(g14851,g12505,g7738);
	nand 	XG4397 	(g14807,g12453,g7738);
	and 	XG4398 	(g14438,g10726,g1087);
	nand 	XG4399 	(g7857,I12242,I12241);
	not 	XG4400 	(g10542,g7196);
	nor 	XG4401 	(g14392,g9537,g12114);
	not 	XG4402 	(g12886,g10393);
	nand 	XG4403 	(g8873,I12850,I12849);
	nand 	XG4404 	(g13273,g10699,g1459);
	nand 	XG4405 	(g13315,g10715,g1459);
	not 	XG4406 	(g11170,g8476);
	not 	XG4407 	(g11512,g7634);
	nand 	XG4408 	(g14407,g9807,g12008);
	not 	XG4409 	(g14545,g12768);
	not 	XG4410 	(g11510,g7633);
	nand 	XG4411 	(g13121,g8411,g11117);
	not 	XG4412 	(g10741,g8411);
	not 	XG4413 	(g10761,g8411);
	nand 	XG4414 	(I14186,I14185,g8442);
	not 	XG4415 	(g11981,I14823);
	or 	XG4416 	(g14030,g11046,g11037);
	nand 	XG4417 	(g9823,I13384,I13383);
	not 	XG4418 	(g12879,g10381);
	not 	XG4419 	(g10504,g8763);
	not 	XG4420 	(g12884,g10392);
	not 	XG4421 	(g10678,I13990);
	not 	XG4422 	(g11192,g8038);
	or 	XG4423 	(g13973,g11028,g11024);
	not 	XG4424 	(g11592,I14537);
	nand 	XG4425 	(I14258,I14257,g8154);
	not 	XG4426 	(I14833,g10142);
	nand 	XG4427 	(g10336,I13751,I13750);
	nand 	XG4428 	(g9904,I13444,I13443);
	or 	XG4429 	(g13570,g11130,g9223);
	and 	XG4430 	(I16143,g11445,g11491,g8751);
	and 	XG4431 	(g14506,g10755,g1430);
	or 	XG4432 	(g13699,g10947,g10921);
	not 	XG4433 	(g14004,g11149);
	not 	XG4434 	(g12107,g9687);
	and 	XG4435 	(g14148,g10632,g884);
	and 	XG4436 	(g14126,g10632,g881);
	nand 	XG4437 	(g14892,g12515,g12700);
	nand 	XG4438 	(g15018,g12515,g12739);
	nand 	XG4439 	(g14858,g12515,g7766);
	nand 	XG4440 	(g12512,g10312,g7766);
	nand 	XG4441 	(g14968,g10312,g12739);
	nand 	XG4442 	(g14810,g10312,g12700);
	and 	XG4443 	(g10869,g5881,g5873,g7766);
	and 	XG4444 	(g14614,g11997,g11975);
	nand 	XG4445 	(I14884,I14883,g9500);
	nor 	XG4446 	(g11771,g4185,g8921);
	not 	XG4447 	(g12944,g12659);
	nand 	XG4448 	(g14895,g12571,g7766);
	nand 	XG4449 	(g14813,g12824,g7766);
	not 	XG4450 	(g12009,I14862);
	nand 	XG4451 	(g13708,g8507,g11200);
	nor 	XG4452 	(g12492,g5164,g5170,g7704);
	nand 	XG4453 	(g14755,g12772,g12593);
	nand 	XG4454 	(g14841,g12443,g12593);
	nand 	XG4455 	(g13134,g8470,g11134);
	nand 	XG4456 	(g14981,g12632,g12785);
	nand 	XG4457 	(g15014,g12680,g12785);
	nor 	XG4458 	(g12716,g6549,g6555,g7812);
	not 	XG4459 	(g10627,I13968);
	nand 	XG4460 	(g13739,g11261,g11773);
	nand 	XG4461 	(g13634,g11261,g11797);
	not 	XG4462 	(g13995,g11261);
	not 	XG4463 	(g10429,g7148);
	not 	XG4464 	(g11249,g8405);
	nand 	XG4465 	(g7887,I12279,I12278);
	not 	XG4466 	(g11724,I14593);
	nor 	XG4467 	(g12067,g7051,g5990);
	nand 	XG4468 	(g12577,g6044,g5990,g7051);
	and 	XG4469 	(g11139,g9935,g5976,g7051,g5990);
	nor 	XG4470 	(g12129,g7051,g9992);
	not 	XG4471 	(g12898,g10405);
	nand 	XG4472 	(I14817,I14816,g9962);
	not 	XG4473 	(g10981,I14119);
	and 	XG4474 	(g13035,g11033,g8497);
	and 	XG4475 	(g13493,g11866,g9880);
	not 	XG4476 	(g12889,g10396);
	not 	XG4477 	(g10533,g8795);
	nand 	XG4478 	(g10738,g10308,g6961);
	nand 	XG4479 	(g9975,I13520,I13519);
	nor 	XG4480 	(g11194,g6875,g3288);
	nand 	XG4481 	(g11479,g3347,g3288,g6875);
	and 	XG4482 	(g10721,g8481,g3274,g6875,g3288);
	nor 	XG4483 	(g11217,g6875,g8531);
	not 	XG4484 	(g12859,g10366);
	nand 	XG4485 	(I15004,I15002,g1700);
	not 	XG4486 	(g12381,I15223);
	nor 	XG4487 	(g12002,g7004,g5297);
	nand 	XG4488 	(g12449,g5352,g5297,g7004);
	and 	XG4489 	(g10588,g5297,g7004);
	and 	XG4490 	(g11111,g9780,g5283,g7004,g5297);
	nor 	XG4491 	(g12059,g7004,g9853);
	not 	XG4492 	(g12890,g10397);
	nand 	XG4493 	(g13432,g10831,g4793);
	nor 	XG4494 	(g14418,g9594,g12151);
	not 	XG4495 	(g12900,g10406);
	and 	XG4496 	(g13523,g12246,g7046);
	nand 	XG4497 	(g13330,g11006,g4664);
	nor 	XG4498 	(g14446,g9644,g12190);
	nand 	XG4499 	(g14170,g11537,g11715);
	nand 	XG4500 	(g14082,g11537,g11697);
	nand 	XG4501 	(g14058,g11537,g7121);
	nand 	XG4502 	(g14142,g8958,g11715);
	nand 	XG4503 	(g14021,g8958,g11697);
	nand 	XG4504 	(g11534,g8958,g7121);
	and 	XG4505 	(g12735,g3881,g3873,g7121);
	nand 	XG4506 	(I14398,g3654,g8542);
	not 	XG4507 	(g14237,g11666);
	nand 	XG4508 	(g14085,g11584,g7121);
	nand 	XG4509 	(g14024,g11763,g7121);
	not 	XG4510 	(g11143,g8032);
	nor 	XG4511 	(g11448,g8790,g4191);
	not 	XG4512 	(g11398,I14409);
	not 	XG4513 	(g10762,g8470);
	not 	XG4514 	(g10794,g8470);
	nand 	XG4515 	(g7223,I11879,I11878);
	not 	XG4516 	(I15033,g10273);
	not 	XG4517 	(g12367,I15205);
	not 	XG4518 	(g12903,g10411);
	nand 	XG4519 	(g9966,I13499,I13498);
	not 	XG4520 	(g12862,g10370);
	nor 	XG4521 	(g14792,g10611,g10618,g10623,g10653);
	and 	XG4522 	(g14644,g10605,g10610);
	not 	XG4523 	(g11467,g7623);
	not 	XG4524 	(g11450,I14455);
	not 	XG4525 	(g11128,g7993);
	not 	XG4526 	(g12867,g10375);
	nand 	XG4527 	(g14999,g12824,g12739);
	nand 	XG4528 	(g14855,g12824,g12700);
	nand 	XG4529 	(g14933,g12571,g12700);
	nand 	XG4530 	(g14735,g12571,g12739);
	nand 	XG4531 	(g14127,g11435,g11653);
	nand 	XG4532 	(g13889,g11435,g11566);
	nand 	XG4533 	(g13892,g11473,g11653);
	nand 	XG4534 	(g13915,g11473,g11566);
	not 	XG4535 	(g14208,g11563);
	and 	XG4536 	(g13048,g11043,g8558);
	nand 	XG4537 	(I14368,g3303,g8481);
	not 	XG4538 	(g12864,g10373);
	nor 	XG4539 	(g11207,g6905,g3639);
	not 	XG4540 	(g12863,g10371);
	nand 	XG4541 	(g11444,g8733,g6918,g6905);
	nor 	XG4542 	(g11238,g6905,g8584);
	not 	XG4543 	(g11519,g8481);
	not 	XG4544 	(g12869,g10376);
	and 	XG4545 	(g13080,g11357,g6923);
	and 	XG4546 	(g11166,I14225,g8296,g269,g8363);
	nand 	XG4547 	(g13795,g401,g11216);
	nor 	XG4548 	(g14816,g12252,g10166);
	or 	XG4549 	(g13794,g10684,g7396);
	not 	XG4550 	(g11640,I14550);
	nor 	XG4551 	(g12645,g6961,g4467);
	nand 	XG4552 	(g12767,g6961,g4467);
	nand 	XG4553 	(g12796,g6961,g4467);
	not 	XG4554 	(I13802,g6971);
	not 	XG4555 	(g10658,I13979);
	and 	XG4556 	(g14586,g11970,g11953);
	not 	XG4557 	(g12896,g10402);
	and 	XG4558 	(g13507,g12198,g7023);
	nor 	XG4559 	(g14212,g10537,g5373);
	nand 	XG4560 	(I15263,I15262,g10081);
	not 	XG4561 	(g11509,g7632);
	and 	XG4562 	(g14202,g10632,g869);
	and 	XG4563 	(g14190,g10632,g859);
	and 	XG4564 	(g14680,g12053,g12024);
	and 	XG4565 	(I16618,g12293,g12341,g10124);
	nand 	XG4566 	(g10041,I13566,I13565);
	nor 	XG4567 	(g14752,g10040,g12540);
	nand 	XG4568 	(g14665,g12798,g12604);
	nand 	XG4569 	(g14959,g12798,g12695);
	nand 	XG4570 	(g14927,g10281,g12695);
	nand 	XG4571 	(g14956,g10281,g12604);
	not 	XG4572 	(g12430,I15250);
	and 	XG4573 	(g14791,g10909,g1146);
	not 	XG4574 	(g13729,g10951);
	not 	XG4575 	(g13595,g10951);
	not 	XG4576 	(g13569,g10951);
	not 	XG4577 	(g13624,g10951);
	nand 	XG4578 	(g14868,g12680,g12755);
	nand 	XG4579 	(g14822,g12632,g12755);
	nand 	XG4580 	(g12915,g12632,g12806);
	nand 	XG4581 	(g14825,g12680,g12806);
	not 	XG4582 	(g12945,g12467);
	nand 	XG4583 	(g14157,g11763,g11715);
	nand 	XG4584 	(g14055,g11763,g11697);
	nand 	XG4585 	(g13963,g11584,g11715);
	nand 	XG4586 	(g14116,g11584,g11697);
	nand 	XG4587 	(I14187,I14185,g3470);
	nand 	XG4588 	(g14918,g12772,g12646);
	nand 	XG4589 	(g14627,g12772,g12553);
	nand 	XG4590 	(g14723,g12772,g7704);
	nand 	XG4591 	(g14800,g12443,g7704);
	nand 	XG4592 	(g14659,g12443,g12646);
	nand 	XG4593 	(g14683,g12443,g12553);
	not 	XG4594 	(g12563,g9864);
	not 	XG4595 	(g13103,g10905);
	not 	XG4596 	(g13215,g10909);
	not 	XG4597 	(g13188,g10909);
	not 	XG4598 	(g13175,g10909);
	not 	XG4599 	(g11147,g8417);
	nand 	XG4600 	(g8238,I12470,I12469);
	nand 	XG4601 	(g14521,g5428,g12170);
	nand 	XG4602 	(g14547,g12201,g9439);
	nand 	XG4603 	(g7598,I12076,I12075);
	nand 	XG4604 	(g12644,g4531,g10233);
	not 	XG4605 	(g12878,g10386);
	not 	XG4606 	(g12882,g10389);
	not 	XG4607 	(I13805,g6976);
	not 	XG4608 	(g10805,I14046);
	not 	XG4609 	(g11183,g8135);
	not 	XG4610 	(g12836,g10351);
	nand 	XG4611 	(I14765,I14764,g9808);
	not 	XG4612 	(g13869,g10831);
	not 	XG4613 	(g13297,g10831);
	not 	XG4614 	(g14231,g12246);
	or 	XG4615 	(g13997,g11036,g11029);
	nand 	XG4616 	(g14573,g12249,g9506);
	nand 	XG4617 	(g9912,I13464,I13463);
	nand 	XG4618 	(I15042,I15041,g9752);
	not 	XG4619 	(I13779,g6868);
	nand 	XG4620 	(g9310,I13079,I13078);
	nand 	XG4621 	(g14741,g10421,g12711);
	nand 	XG4622 	(g14817,g12622,g12711);
	not 	XG4623 	(I14800,g10107);
	nand 	XG4624 	(I14482,I14480,g655);
	not 	XG4625 	(g12870,g10374);
	not 	XG4626 	(g11471,g7626);
	not 	XG4627 	(g11576,g8542);
	nand 	XG4628 	(g14333,g11892,g11990,g12014,g12042);
	nand 	XG4629 	(g12910,g10601,g11002);
	not 	XG4630 	(g10804,g9772);
	nand 	XG4631 	(g13870,g4732,g11773);
	nor 	XG4632 	(g14872,g12364,g6736);
	nand 	XG4633 	(g12686,g6736,g6682,g7097);
	nand 	XG4634 	(g13855,g11804,g4944);
	and 	XG4635 	(g13384,g11804,g4944);
	not 	XG4636 	(g12888,g10395);
	not 	XG4637 	(g14215,g12198);
	nand 	XG4638 	(g7201,I11866,I11865);
	nand 	XG4639 	(I14205,I14204,g8508);
	nand 	XG4640 	(g9528,I13184,I13183);
	nand 	XG4641 	(I14259,I14257,g3133);
	not 	XG4642 	(g12860,g10368);
	not 	XG4643 	(g12841,g10357);
	not 	XG4644 	(g13521,g11357);
	or 	XG4645 	(g13300,g10676,g10656);
	nand 	XG4646 	(g13851,g11360,g8224);
	nand 	XG4647 	(I15175,I15174,g9977);
	nor 	XG4648 	(g14793,g12228,g2988);
	nor 	XG4649 	(g14754,g2988,g12821);
	not 	XG4650 	(g12907,g10415);
	nand 	XG4651 	(g7897,I12289,I12288);
	nand 	XG4652 	(g13886,g4922,g11804);
	not 	XG4653 	(g10532,g10233);
	not 	XG4654 	(g10620,g10233);
	not 	XG4655 	(g10509,g10233);
	not 	XG4656 	(g10606,g10233);
	not 	XG4657 	(g10607,g10233);
	not 	XG4658 	(I14192,g10233);
	not 	XG4659 	(I14346,g10233);
	not 	XG4660 	(g10487,g10233);
	not 	XG4661 	(g10597,g10233);
	not 	XG4662 	(g10572,g10233);
	not 	XG4663 	(g10612,g10233);
	not 	XG4664 	(g10613,g10233);
	not 	XG4665 	(g12820,g10233);
	not 	XG4666 	(g10571,g10233);
	nor 	XG4667 	(g14713,g9974,g12483);
	not 	XG4668 	(g11428,g7615);
	nor 	XG4669 	(g14772,g12252,g6044);
	nand 	XG4670 	(g12462,g10190,g7064,g7051);
	not 	XG4671 	(g12930,g12347);
	not 	XG4672 	(g13120,g10632);
	not 	XG4673 	(g13140,g10632);
	not 	XG4674 	(g13173,g10632);
	not 	XG4675 	(g13239,g10632);
	not 	XG4676 	(g13255,g10632);
	not 	XG4677 	(g13132,g10632);
	not 	XG4678 	(g13209,g10632);
	not 	XG4679 	(g13142,g10632);
	nand 	XG4680 	(g13176,g1404,g1322,g7675,g10715);
	nand 	XG4681 	(g13137,g1404,g1322,g7675,g10699);
	not 	XG4682 	(g10417,g7117);
	nor 	XG4683 	(g12026,g9340,g9417);
	not 	XG4684 	(g12487,g9340);
	not 	XG4685 	(I14602,g9340);
	not 	XG4686 	(I14650,g9340);
	not 	XG4687 	(I14690,g9340);
	not 	XG4688 	(g12337,g9340);
	not 	XG4689 	(I14633,g9340);
	not 	XG4690 	(I15831,g10416);
	not 	XG4691 	(I16917,g10582);
	not 	XG4692 	(g11402,g7594);
	not 	XG4693 	(g12845,g10358);
	not 	XG4694 	(g12842,g10355);
	nand 	XG4695 	(g13102,g10759,g7523);
	not 	XG4696 	(g10816,I14054);
	nor 	XG4697 	(g13501,g11881,g3368);
	not 	XG4698 	(g10815,g9917);
	not 	XG4699 	(g12872,g10379);
	nand 	XG4700 	(I15342,I15340,g2541);
	and 	XG4701 	(g14567,g10552,g10568);
	or 	XG4702 	(g13289,g10624,g10619);
	nand 	XG4703 	(g9908,I13454,I13453);
	not 	XG4704 	(g14209,g11415);
	not 	XG4705 	(g14405,g12170);
	not 	XG4706 	(g11325,g7543);
	not 	XG4707 	(g11498,I14475);
	and 	XG4708 	(g14643,g12023,g11998);
	not 	XG4709 	(g12760,g10272);
	nand 	XG4710 	(I14611,I14609,g8678);
	not 	XG4711 	(g11048,I14158);
	nand 	XG4712 	(I14352,I14350,g8848);
	not 	XG4713 	(g13504,g11303);
	or 	XG4714 	(g13295,g10655,g10625);
	not 	XG4715 	(g14186,g11346);
	not 	XG4716 	(g12874,g10383);
	nor 	XG4717 	(g14914,g12797,g12822);
	not 	XG4718 	(g11371,g7565);
	and 	XG4719 	(g13632,g12228,g10232);
	not 	XG4720 	(g14432,g12311);
	not 	XG4721 	(g13663,g10971);
	not 	XG4722 	(g13596,g10971);
	not 	XG4723 	(g13763,g10971);
	not 	XG4724 	(g13625,g10971);
	nand 	XG4725 	(g8359,I12546,I12545);
	nand 	XG4726 	(g13797,g11273,g8102);
	not 	XG4727 	(g11367,I14381);
	not 	XG4728 	(I15295,g8515);
	not 	XG4729 	(g11164,g8085);
	not 	XG4730 	(g12705,g7051);
	nand 	XG4731 	(g12972,g10578,g7209);
	nand 	XG4732 	(g11410,g8696,g6895,g6875);
	not 	XG4733 	(g11468,g7624);
	not 	XG4734 	(I14708,g9417);
	not 	XG4735 	(g12378,g9417);
	not 	XG4736 	(g12543,g9417);
	not 	XG4737 	(I14653,g9417);
	not 	XG4738 	(g12598,g7004);
	or 	XG4739 	(g13972,g11203,g11232);
	nand 	XG4740 	(g13779,g11283,g11804);
	nand 	XG4741 	(g13676,g11283,g11834);
	not 	XG4742 	(g14029,g11283);
	or 	XG4743 	(g13914,g11380,g8643);
	not 	XG4744 	(g12818,g8792);
	not 	XG4745 	(I14579,g8792);
	not 	XG4746 	(I14623,g8925);
	not 	XG4747 	(g10531,g8925);
	not 	XG4748 	(g10503,g8879);
	not 	XG4749 	(g10419,g8821);
	not 	XG4750 	(g12868,g10377);
	nand 	XG4751 	(g13217,g10808,g4082);
	and 	XG4752 	(g13063,g10808,g8567);
	not 	XG4753 	(g11560,g7647);
	nor 	XG4754 	(g14413,g9638,g11914);
	not 	XG4755 	(g12640,I15382);
	not 	XG4756 	(g11608,g7659);
	not 	XG4757 	(g11403,g7595);
	nor 	XG4758 	(g12137,g7097,g6682);
	not 	XG4759 	(g12906,g10413);
	nand 	XG4760 	(g12590,g10229,g7110,g7097);
	nor 	XG4761 	(g12211,g7097,g10099);
	not 	XG4762 	(g14503,g12256);
	nand 	XG4763 	(I15254,I15253,g10078);
	nand 	XG4764 	(g14489,g5084,g12126);
	nand 	XG4765 	(g14520,g12163,g9369);
	and 	XG4766 	(g14615,g10587,g10604);
	or 	XG4767 	(g13296,g10657,g10626);
	nor 	XG4768 	(g13939,g11173,g8822,g4899);
	nor 	XG4769 	(g13910,g11173,g4975,g4899);
	nand 	XG4770 	(g12155,g7717,g7753);
	not 	XG4771 	(I14668,g7753);
	not 	XG4772 	(I14687,g7753);
	not 	XG4773 	(I14727,g7753);
	not 	XG4774 	(I14761,g7753);
	and 	XG4775 	(g11032,g7717,g9354);
	not 	XG4776 	(g11373,g7566);
	nand 	XG4777 	(g14993,g12453,g12695);
	nand 	XG4778 	(g14688,g12453,g12604);
	nand 	XG4779 	(g14691,g12505,g12695);
	nand 	XG4780 	(g14727,g12505,g12604);
	not 	XG4781 	(g12936,g12601);
	nand 	XG4782 	(g14434,g11945,g6415);
	nand 	XG4783 	(g14899,g10421,g12744);
	nand 	XG4784 	(g15024,g10421,g12780);
	nand 	XG4785 	(g14974,g12622,g12744);
	nand 	XG4786 	(g14776,g12622,g12780);
	not 	XG4787 	(g12834,g10349);
	nand 	XG4788 	(g7869,I12253,I12252);
	nand 	XG4789 	(g13871,g11834,g4955);
	and 	XG4790 	(g13411,g11834,g4955);
	not 	XG4791 	(g12880,g10387);
	nor 	XG4792 	(g14416,g9541,g12148);
	not 	XG4793 	(g12937,g12419);
	nand 	XG4794 	(g9258,I13045,I13044);
	or 	XG4795 	(g13095,g1287,g11374);
	not 	XG4796 	(I13872,g7474);
	not 	XG4797 	(I14660,g9746);
	not 	XG4798 	(g12790,g7097);
	not 	XG4799 	(g11404,g7596);
	nand 	XG4800 	(I14277,I14275,g3484);
	not 	XG4801 	(g12922,g12297);
	not 	XG4802 	(g11868,g9185);
	not 	XG4803 	(I14630,g7717);
	not 	XG4804 	(I14705,g7717);
	not 	XG4805 	(I14730,g7717);
	not 	XG4806 	(I14647,g7717);
	not 	XG4807 	(I14702,g7717);
	not 	XG4808 	(I14684,g7717);
	not 	XG4809 	(I14644,g7717);
	not 	XG4810 	(I14671,g7717);
	not 	XG4811 	(g11819,g7717);
	nand 	XG4812 	(g12491,g6961,g4462,g7285);
	nand 	XG4813 	(g12819,g6961,g9848);
	nand 	XG4814 	(g10737,g9848,g6961);
	not 	XG4815 	(g11652,g7674);
	nand 	XG4816 	(g14601,g6466,g12318);
	or 	XG4817 	(g14062,g11116,g11047);
	nand 	XG4818 	(g14638,g12361,g9626);
	not 	XG4819 	(g14504,g12361);
	nand 	XG4820 	(g9825,I13392,I13391);
	not 	XG4821 	(g14251,g12308);
	nand 	XG4822 	(g13346,g11012,g4854);
	nand 	XG4823 	(I14248,I14247,g1322);
	not 	XG4824 	(g12844,g10360);
	and 	XG4825 	(g14588,g11974,g11957);
	not 	XG4826 	(g11290,I14326);
	and 	XG4827 	(g14613,g10585,g10602);
	not 	XG4828 	(g12672,g10003);
	not 	XG4829 	(g12893,g10391);
	not 	XG4830 	(g11234,g8355);
	nand 	XG4831 	(I14885,I14883,g5489);
	not 	XG4832 	(g12837,g10354);
	not 	XG4833 	(g11709,I14584);
	nor 	XG4834 	(g14515,g9761,g12225);
	nor 	XG4835 	(g14395,g9542,g12118);
	nand 	XG4836 	(g8737,I12730,I12729);
	not 	XG4837 	(g13301,g10862);
	not 	XG4838 	(g13885,g10862);
	not 	XG4839 	(g13594,g11012);
	nor 	XG4840 	(g14364,g9415,g12083);
	not 	XG4841 	(I14749,g10031);
	not 	XG4842 	(I14830,g10141);
	nand 	XG4843 	(g9830,I13403,I13402);
	and 	XG4844 	(g14537,g10529,g10550);
	nor 	XG4845 	(g14272,g10598,g6411);
	not 	XG4846 	(g13976,g11130);
	not 	XG4847 	(I14899,g10198);
	and 	XG4848 	(g14565,g11952,g11934);
	nand 	XG4849 	(g12629,g7142,g7812);
	nand 	XG4850 	(g14908,g10491,g7812);
	and 	XG4851 	(g10887,g6573,g6565,g7812);
	and 	XG4852 	(g14641,g12020,g11994);
	nand 	XG4853 	(I15255,I15253,g1848);
	not 	XG4854 	(g12861,g10367);
	and 	XG4855 	(g13046,g11270,g6870);
	not 	XG4856 	(g12892,g10398);
	and 	XG4857 	(g13491,g12160,g6999);
	not 	XG4858 	(I14663,g9747);
	not 	XG4859 	(g11686,I14567);
	not 	XG4860 	(g10530,g8922);
	not 	XG4861 	(I14589,g8818);
	not 	XG4862 	(g10418,g8818);
	not 	XG4863 	(g11324,g7542);
	nor 	XG4864 	(g13378,g11017,g11374);
	not 	XG4865 	(g12929,g12550);
	not 	XG4866 	(I16010,g11148);
	not 	XG4867 	(g12811,g10319);
	not 	XG4868 	(g14535,g12318);
	not 	XG4869 	(g14342,g12163);
	not 	XG4870 	(g14376,g12126);
	not 	XG4871 	(I16898,g10615);
	nand 	XG4872 	(g7885,I12271,I12270);
	not 	XG4873 	(g12840,g10356);
	nand 	XG4874 	(g14950,g12632,g7812);
	nand 	XG4875 	(g14984,g12680,g7812);
	nand 	XG4876 	(I14992,I14991,g9685);
	not 	XG4877 	(g13483,g11270);
	not 	XG4878 	(g13141,g11374);
	nor 	XG4879 	(g14751,g10603,g10609,g10617,g10622);
	nor 	XG4880 	(g14449,g9653,g12194);
	not 	XG4881 	(g10554,g8974);
	not 	XG4882 	(g10475,g8844);
	not 	XG4883 	(g13715,g10573);
	not 	XG4884 	(g13679,g10573);
	not 	XG4885 	(g13621,g10573);
	not 	XG4886 	(g13655,g10573);
	not 	XG4887 	(g11930,g9281);
	not 	XG4888 	(g14275,g12358);
	not 	XG4889 	(g13637,g10556);
	not 	XG4890 	(g13675,g10556);
	not 	XG4891 	(g13620,g10556);
	not 	XG4892 	(g13593,g10556);
	not 	XG4893 	(g11431,g7618);
	not 	XG4894 	(g11202,I14267);
	not 	XG4895 	(g12895,g10403);
	not 	XG4896 	(g12921,g12228);
	not 	XG4897 	(g14197,g12160);
	not 	XG4898 	(g10498,g7161);
	not 	XG4899 	(g10812,I14050);
	nand 	XG4900 	(g8913,I12878,I12877);
	not 	XG4901 	(g11547,I14505);
	not 	XG4902 	(I15800,g11607);
	nand 	XG4903 	(I14351,I14350,g8890);
	not 	XG4904 	(g11268,g7515);
	not 	XG4905 	(g13133,g11330);
	nand 	XG4906 	(I15043,I15041,g1834);
	not 	XG4907 	(g12656,g7028);
	nand 	XG4908 	(g9750,I13336,I13335);
	nand 	XG4909 	(I15129,I15128,g9914);
	not 	XG4910 	(I15316,g10087);
	not 	XG4911 	(g10830,g10087);
	not 	XG4912 	(g12975,g12752);
	nand 	XG4913 	(I14993,I14991,g6527);
	not 	XG4914 	(g12894,g10401);
	not 	XG4915 	(I14745,g10029);
	not 	XG4916 	(g12914,g12235);
	not 	XG4917 	(g12881,g10388);
	not 	XG4918 	(g11663,g6905);
	not 	XG4919 	(g12614,g9935);
	not 	XG4920 	(g11215,g8285);
	not 	XG4921 	(g14406,g12249);
	not 	XG4922 	(g11425,g7640);
	not 	XG4923 	(g11615,g6875);
	not 	XG4924 	(g13506,g10808);
	not 	XG4925 	(g14377,g12201);
	nand 	XG4926 	(I15176,I15174,g2661);
	not 	XG4927 	(I16024,g11171);
	not 	XG4928 	(g13565,g11006);
	not 	XG4929 	(g10570,g9021);
	not 	XG4930 	(g13626,g11273);
	not 	XG4931 	(g10502,g8876);
	not 	XG4932 	(g13026,g11018);
	not 	XG4933 	(g10474,g8841);
	not 	XG4934 	(I14576,g8791);
	not 	XG4935 	(g13707,g11360);
	not 	XG4936 	(g10776,I14033);
	not 	XG4937 	(g10685,I13995);
	not 	XG4938 	(g14226,g11618);
	not 	XG4939 	(I13759,g6754);
	not 	XG4940 	(I13762,g6755);
	not 	XG4941 	(g12873,g10380);
	not 	XG4942 	(I14016,g9104);
	not 	XG4943 	(I14069,g9104);
	not 	XG4944 	(I14006,g9104);
	not 	XG4945 	(I16231,g10520);
	not 	XG4946 	(g12793,g10287);
	not 	XG4947 	(I14305,g8805);
	not 	XG4948 	(g10857,g8712);
	nor 	XG4949 	(g14393,g9488,g12115);
	or 	XG4950 	(g12911,g12768,g10278);
	nand 	XG4951 	(g12414,g10165,g7041,g7028);
	nor 	XG4952 	(g14731,g12204,g5698);
	nor 	XG4953 	(g14726,g12166,g10090);
	nand 	XG4954 	(I14854,I14853,g9433);
	nand 	XG4955 	(I15130,I15128,g2527);
	nor 	XG4956 	(g14394,g9414,g12116);
	nand 	XG4957 	(I14610,I14609,g8993);
	nand 	XG4958 	(g14378,g9731,g11979);
	nand 	XG4959 	(g14146,g691,g11020);
	nand 	XG4960 	(g13945,g11740,g691);
	nand 	XG4961 	(I14290,I14289,g8282);
	nor 	XG4962 	(g14568,g9915,g12000);
	nand 	XG4963 	(g13266,g9843,g9920,g12440);
	nand 	XG4964 	(g13248,g9843,g12399,g9985);
	nand 	XG4965 	(g13283,g9843,g12399,g12440);
	nand 	XG4966 	(g12971,g10664,g8977,g9024);
	nand 	XG4967 	(I14714,I14712,g5128);
	nand 	XG4968 	(I15299,I15298,g10112);
	nand 	XG4969 	(I14517,I14516,g10147);
	nor 	XG4970 	(g14367,g12289,g9547);
	nor 	XG4971 	(g14339,g2735,g12289);
	and 	XG4972 	(g13038,g11034,g8509);
	nand 	XG4973 	(I14206,I14204,g3821);
	nand 	XG4974 	(I14170,I14169,g8389);
	nand 	XG4975 	(g13513,g8002,g11815,g1351);
	nand 	XG4976 	(I14924,I14923,g9558);
	nor 	XG4977 	(g14642,g9829,g12374);
	and 	XG4978 	(g13524,g11910,g9995);
	or 	XG4979 	(g13077,g943,g11330);
	or 	XG4980 	(g13597,g11149,g9247);
	nand 	XG4981 	(I14766,I14764,g5821);
	nand 	XG4982 	(g13850,g8396,g11279);
	nand 	XG4983 	(g14600,g12311,g9564);
	nand 	XG4984 	(g14574,g6120,g12256);
	nand 	XG4985 	(g12342,g10129,g7018,g7004);
	nor 	XG4986 	(g14687,g12166,g5352);
	nor 	XG4987 	(g12093,g7028,g9924);
	nand 	XG4988 	(g12511,g5698,g5644,g7028);
	nor 	XG4989 	(g12029,g7028,g5644);
	nor 	XG4990 	(g14611,g9749,g12333);
	nand 	XG4991 	(g14505,g9961,g12073);
	nand 	XG4992 	(I15307,I15306,g10116);
	and 	XG4993 	(g14585,g10905,g1141);
	nand 	XG4994 	(I15364,I15363,g10182);
	nand 	XG4995 	(I15335,I15333,g2116);
	nor 	XG4996 	(g14396,g9489,g12119);
	not 	XG4997 	(g13706,g11280);
	nor 	XG4998 	(g14538,g9828,g11973);
	nor 	XG4999 	(g14121,g12259,g8891);
	nor 	XG5000 	(g14337,g9284,g12049);
	nand 	XG5001 	(I15213,I15212,g10035);
	and 	XG5002 	(g13436,g11811,g9721);
	nand 	XG5003 	(I14734,I14733,g9732);
	nor 	XG5004 	(g13989,g11309,g8697);
	nand 	XG5005 	(I14855,I14853,g5142);
	nor 	XG5006 	(g14003,g11083,g9003);
	nor 	XG5007 	(g13996,g11173,g8822,g8938);
	nor 	XG5008 	(g13971,g11173,g4975,g8938);
	nand 	XG5009 	(g14089,g4717,g11755);
	nand 	XG5010 	(g14317,g11862,g5033);
	nand 	XG5011 	(g12524,g10212,g7087,g7074);
	nor 	XG5012 	(g14821,g12314,g6390);
	nand 	XG5013 	(I15300,I15298,g1982);
	and 	XG5014 	(g13525,g11911,g10019);
	nor 	XG5015 	(g14360,g9484,g12078);
	nor 	XG5016 	(g14767,g12204,g10130);
	nand 	XG5017 	(I14509,I14508,g370);
	nand 	XG5018 	(g13884,g4727,g11797);
	and 	XG5019 	(g13025,g11026,g8431);
	and 	XG5020 	(I16111,g11381,g11409,g8691);
	or 	XG5021 	(g13091,g10796,g319,g329);
	nor 	XG5022 	(g11185,g6804,g8183,g8038);
	or 	XG5023 	(g13660,g12527,g8183);
	or 	XG5024 	(g13623,g12527,g482);
	nor 	XG5025 	(g14444,g9692,g11936);
	nor 	XG5026 	(g14447,g9698,g11938);
	nand 	XG5027 	(g10754,g8411,g7913,g7936);
	nand 	XG5028 	(g14344,g11885,g5377);
	nor 	XG5029 	(g14911,g12364,g10213);
	nor 	XG5030 	(g14712,g9971,g12479);
	nor 	XG5031 	(g14450,g9598,g12195);
	and 	XG5032 	(g14831,g10909,g1152);
	nor 	XG5033 	(g14033,g12259,g8808);
	nand 	XG5034 	(I15122,I15121,g9910);
	nor 	XG5035 	(g14513,g9754,g12222);
	nand 	XG5036 	(g15042,g10491,g12806);
	nand 	XG5037 	(g14947,g10491,g12785);
	nand 	XG5038 	(g14782,g10491,g12755);
	nand 	XG5039 	(g15033,g7142,g12806);
	nand 	XG5040 	(g14905,g7142,g12785);
	nand 	XG5041 	(g15039,g7142,g12755);
	nand 	XG5042 	(g14546,g9613,g12125);
	nand 	XG5043 	(g12933,g10515,g7150);
	nor 	XG5044 	(g14391,g9585,g12112);
	and 	XG5045 	(g13287,g11472,g1221);
	nand 	XG5046 	(g14433,g9890,g12035);
	nand 	XG5047 	(g11405,g2748,g6856,g2735,g2741);
	nor 	XG5048 	(g12123,g2748,g6856);
	nor 	XG5049 	(g12377,g9708,g2748,g6856);
	nand 	XG5050 	(g10775,g8470,g7943,g7960);
	and 	XG5051 	(g13383,g11797,g4765);
	nand 	XG5052 	(g13854,g11797,g4765);
	and 	XG5053 	(g13542,g11927,g10053);
	nand 	XG5054 	(I14957,I14955,g6181);
	and 	XG5055 	(g14180,g10632,g872);
	and 	XG5056 	(g10476,I13862,g7259,g7244);
	nand 	XG5057 	(g13495,g7972,g11786,g1008);
	and 	XG5058 	(g13509,g11889,g9951);
	nor 	XG5059 	(g14640,g9824,g12371);
	nor 	XG5060 	(g14362,g9338,g12080);
	nor 	XG5061 	(g14445,g9693,g12188);
	nor 	XG5062 	(g14176,g12259,g9044);
	nor 	XG5063 	(g14516,g9704,g12227);
	nor 	XG5064 	(g14539,g9833,g11977);
	nor 	XG5065 	(g13947,g11083,g8948);
	nor 	XG5066 	(g14397,g9416,g12120);
	and 	XG5067 	(g10590,I13937,g7392,g7246);
	nand 	XG5068 	(I15079,I15078,g9827);
	nand 	XG5069 	(I15052,I15051,g9759);
	nand 	XG5070 	(I14789,I14788,g9891);
	nor 	XG5071 	(g14092,g11083,g8774);
	nor 	XG5072 	(g13970,g11155,g8796,g8883);
	nor 	XG5073 	(g13937,g11155,g4785,g8883);
	nand 	XG5074 	(g13712,g11283,g8984);
	nand 	XG5075 	(g13742,g11283,g11780);
	nor 	XG5076 	(g14540,g9834,g12287);
	nand 	XG5077 	(I15123,I15121,g2102);
	nor 	XG5078 	(g14419,g9546,g12152);
	nor 	XG5079 	(g14036,g11083,g8725);
	nor 	XG5080 	(g14001,g11083,g739);
	nand 	XG5081 	(I14735,I14733,g5475);
	nor 	XG5082 	(g14122,g12259,g8895);
	nor 	XG5083 	(g13512,g12527,g9077);
	nor 	XG5084 	(g13796,g12527,g9158);
	nor 	XG5085 	(g13568,g12527,g8046);
	or 	XG5086 	(g13728,g12527,g6804);
	or 	XG5087 	(g13820,g12527,g9187,g11184);
	nor 	XG5088 	(g14163,g12259,g8997);
	or 	XG5089 	(g12925,g10511,g8928);
	nor 	XG5090 	(g13852,g8347,g11320);
	nor 	XG5091 	(g13202,g10511,g8347);
	nor 	XG5092 	(g13908,g11155,g8796,g4709);
	nand 	XG5093 	(g13672,g11261,g8933);
	nor 	XG5094 	(g13883,g11155,g4785,g4709);
	nand 	XG5095 	(g13709,g11261,g11755);
	nor 	XG5096 	(g14181,g12259,g9083);
	nor 	XG5097 	(g13919,g11276,g3347);
	nand 	XG5098 	(g14637,g9815,g12255);
	nand 	XG5099 	(I15264,I15262,g2273);
	nand 	XG5100 	(g13764,g3072,g11252);
	and 	XG5101 	(g14832,g10939,g1489);
	nor 	XG5102 	(g14091,g12259,g8854);
	nand 	XG5103 	(I15287,g6697,g10061);
	and 	XG5104 	(I16721,g12525,g12589,g10224);
	nand 	XG5105 	(g13666,g8441,g11190);
	nor 	XG5106 	(g14679,g9911,g12437);
	nand 	XG5107 	(g13822,g11306,g8160);
	not 	XG5108 	(I15937,g11676);
	nor 	XG5109 	(g14334,g9337,g12044);
	not 	XG5110 	(I16747,g12729);
	nand 	XG5111 	(I14230,I14228,g8055);
	nor 	XG5112 	(g14037,g11083,g8748);
	nor 	XG5113 	(g14678,g9907,g12432);
	nor 	XG5114 	(g11626,g3857,g3863,g7121);
	nand 	XG5115 	(g13990,g11584,g11669);
	nand 	XG5116 	(g13960,g11537,g11669);
	nand 	XG5117 	(g13929,g11763,g11669);
	nand 	XG5118 	(g14154,g8958,g11669);
	and 	XG5119 	(g14168,g10632,g887);
	or 	XG5120 	(g13385,g9479,g11967);
	nand 	XG5121 	(I14818,I14816,g6513);
	nor 	XG5122 	(g14064,g12259,g9214);
	nand 	XG5123 	(g13667,g11119,g3723);
	nand 	XG5124 	(g13105,g1404,g1322,g7675,g10671);
	nand 	XG5125 	(I13852,I13850,g7397);
	nand 	XG5126 	(g14675,g9898,g12317);
	nor 	XG5127 	(g14707,g12259,g10143);
	nand 	XG5128 	(g13600,g11039,g3021);
	nand 	XG5129 	(g14697,g12824,g12662);
	nand 	XG5130 	(g14768,g12571,g12662);
	nand 	XG5131 	(g14996,g10312,g12662);
	nand 	XG5132 	(g14732,g12515,g12662);
	nor 	XG5133 	(g12609,g5857,g5863,g7766);
	and 	XG5134 	(g14610,g10935,g1484);
	and 	XG5135 	(g13324,g11326,g854);
	nand 	XG5136 	(g13940,g8829,g11707,g8889,g11426);
	nand 	XG5137 	(g14626,g9715,g12159,g9852,g12232);
	nand 	XG5138 	(g13823,g3774,g11313);
	nand 	XG5139 	(g13143,g1061,g979,g7661,g10695);
	nand 	XG5140 	(g13124,g1061,g979,g7661,g10666);
	nand 	XG5141 	(g13093,g1061,g979,g7661,g10649);
	nand 	XG5142 	(I14229,I14228,g979);
	and 	XG5143 	(g13473,g11841,g9797);
	nand 	XG5144 	(g14379,g11907,g5723);
	nand 	XG5145 	(g13284,g1157,g10695);
	nand 	XG5146 	(I13851,I13850,g862);
	and 	XG5147 	(g13060,g11110,g8587);
	nor 	XG5148 	(g14093,g11083,g8833);
	and 	XG5149 	(g14708,g12369,g74);
	nand 	XG5150 	(g14773,g12581,g12711);
	nand 	XG5151 	(g15021,g10341,g12711);
	nor 	XG5152 	(g12667,g6203,g6209,g7791);
	nand 	XG5153 	(g14548,g5774,g12208);
	nand 	XG5154 	(g14572,g9678,g12169);
	nor 	XG5155 	(g14448,g9699,g12192);
	or 	XG5156 	(g12954,g9906,g12186);
	nand 	XG5157 	(g13307,g10695,g1116);
	nand 	XG5158 	(g13846,g10649,g1116);
	nand 	XG5159 	(g13260,g10666,g1116);
	and 	XG5160 	(g13508,g11888,g9927);
	and 	XG5161 	(g10838,g5535,g5527,g7738);
	nand 	XG5162 	(g12450,g10281,g7738);
	nand 	XG5163 	(g14761,g10281,g12651);
	nand 	XG5164 	(g14764,g12798,g7738);
	nand 	XG5165 	(g14804,g12798,g12651);
	nand 	XG5166 	(I14518,I14516,g661);
	nand 	XG5167 	(I15089,I15087,g2393);
	nor 	XG5168 	(g13944,g12259,g10262);
	nor 	XG5169 	(g14414,g9639,g12145);
	not 	XG5170 	(g13736,g11313);
	nand 	XG5171 	(g14343,g9670,g11961);
	and 	XG5172 	(g13047,g11042,g8534);
	nand 	XG5173 	(g11492,g8756,g6941,g6928);
	nor 	XG5174 	(g11255,g6928,g8623);
	and 	XG5175 	(g10756,g8595,g3976,g6928,g3990);
	nor 	XG5176 	(g11225,g6928,g3990);
	not 	XG5177 	(g13665,g11306);
	nor 	XG5178 	(g14000,g12259,g8766);
	nor 	XG5179 	(g14512,g9753,g11955);
	and 	XG5180 	(g12924,g10980,g1570);
	nand 	XG5181 	(g13867,g8449,g11312);
	nand 	XG5182 	(g14258,g11903,g9203);
	nor 	XG5183 	(g13518,g11903,g3719);
	nor 	XG5184 	(g14514,g9760,g11959);
	not 	XG5185 	(g14431,g12208);
	nor 	XG5186 	(g14194,g10515,g5029);
	nor 	XG5187 	(g14027,g11363,g8734);
	nand 	XG5188 	(g14797,g12405,g12593);
	nand 	XG5189 	(g14720,g10266,g12593);
	nand 	XG5190 	(I14427,g4005,g8595);
	nand 	XG5191 	(g14599,g9739,g12207);
	nand 	XG5192 	(g12947,g10561,g7184);
	nor 	XG5193 	(g14228,g10561,g5719);
	and 	XG5194 	(g13294,g11513,g1564);
	nand 	XG5195 	(g11590,g4049,g3990,g6928);
	nor 	XG5196 	(g13994,g11363,g4049);
	and 	XG5197 	(g12920,g10960,g1227);
	nor 	XG5198 	(g14164,g12259,g9000);
	nor 	XG5199 	(g14253,g9217,g12259,g10032);
	nor 	XG5200 	(g13946,g11083,g8651);
	not 	XG5201 	(g13246,g10939);
	not 	XG5202 	(g13216,g10939);
	not 	XG5203 	(g13190,g10939);
	nor 	XG5204 	(g13342,g10935,g10961);
	not 	XG5205 	(g13116,g10935);
	nor 	XG5206 	(g14365,g9339,g12084);
	and 	XG5207 	(g11890,g9155,g7499);
	or 	XG5208 	(g13657,g10616,g7251);
	nand 	XG5209 	(I14291,I14289,g3835);
	and 	XG5210 	(g12641,g3179,g3171,g10295);
	nand 	XG5211 	(g11432,g8864,g10295);
	nand 	XG5212 	(g13948,g8864,g11610);
	nand 	XG5213 	(g13951,g11729,g10295);
	nand 	XG5214 	(g13977,g11729,g11610);
	not 	XG5215 	(g14095,g11326);
	nand 	XG5216 	(g13821,g8340,g11251);
	nand 	XG5217 	(g14223,g11858,g9092);
	and 	XG5218 	(g13247,g11316,g8964);
	or 	XG5219 	(g12981,g9967,g12219);
	nand 	XG5220 	(g14130,g8906,g11621);
	nand 	XG5221 	(g14110,g8906,g11692);
	nand 	XG5222 	(g13983,g8906,g11658);
	nand 	XG5223 	(g13898,g11747,g11621);
	nand 	XG5224 	(g14133,g11747,g11692);
	nand 	XG5225 	(g14015,g11747,g11658);
	nor 	XG5226 	(g14420,g9490,g12153);
	nand 	XG5227 	(I15105,g5313,g9780);
	nor 	XG5228 	(g14090,g12259,g8851);
	nor 	XG5229 	(g14188,g12259,g9162);
	nor 	XG5230 	(g14145,g12259,g8945);
	nor 	XG5231 	(g14278,g9217,g12259,g562);
	and 	XG5232 	(I16129,g11411,g11443,g8728);
	or 	XG5233 	(g13938,g11191,g11213);
	not 	XG5234 	(g13664,g11252);
	nand 	XG5235 	(I15080,I15078,g1968);
	nand 	XG5236 	(g14279,g9246,g12111);
	nor 	XG5237 	(g13480,g11858,g3017);
	nand 	XG5238 	(I15214,I15212,g1714);
	or 	XG5239 	(g13761,g12527,g490);
	nand 	XG5240 	(g14682,g11780,g4933);
	and 	XG5241 	(g13349,g11780,g4933);
	nand 	XG5242 	(g13281,g1099,g10916);
	and 	XG5243 	(g14875,g10939,g1495);
	and 	XG5244 	(g14913,g10939,g1442);
	nand 	XG5245 	(I14925,I14923,g5835);
	nand 	XG5246 	(I15053,I15051,g2259);
	nand 	XG5247 	(g13861,g10671,g1459);
	and 	XG5248 	(g11144,I14198,g246,g8136,g239);
	nand 	XG5249 	(I14790,I14788,g6167);
	nand 	XG5250 	(g14655,g11755,g4743);
	and 	XG5251 	(g13333,g11755,g4743);
	or 	XG5252 	(g13762,g12527,g499);
	nand 	XG5253 	(g13798,g3423,g11280);
	nand 	XG5254 	(g14120,g4907,g11780);
	nand 	XG5255 	(I15365,I15363,g2675);
	nand 	XG5256 	(I15308,I15306,g2407);
	nand 	XG5257 	(I14171,I14169,g3119);
	not 	XG5258 	(g13835,I16150);
	not 	XG5259 	(g14366,I16526);
	not 	XG5260 	(g13680,I16077);
	not 	XG5261 	(g13745,I16102);
	not 	XG5262 	(g12932,I15550);
	not 	XG5263 	(g14338,I16502);
	not 	XG5264 	(g13144,I15773);
	not 	XG5265 	(g14315,I16479);
	not 	XG5266 	(g13782,I16117);
	not 	XG5267 	(g12983,I15600);
	not 	XG5268 	(g13605,I16040);
	not 	XG5269 	(g13416,I15929);
	not 	XG5270 	(g13716,I16090);
	not 	XG5271 	(g13638,I16057);
	not 	XG5272 	(g14336,I16498);
	not 	XG5273 	(g14591,I16709);
	not 	XG5274 	(g14290,I16460);
	not 	XG5275 	(g13329,I15893);
	not 	XG5276 	(g13394,I15915);
	not 	XG5277 	(g13177,I15782);
	not 	XG5278 	(g14314,I16476);
	not 	XG5279 	(g14398,I16555);
	not 	XG5280 	(g12955,I15577);
	not 	XG5281 	(g13350,I15906);
	not 	XG5282 	(g13809,I16135);
	not 	XG5283 	(g14454,I16613);
	not 	XG5284 	(g13191,I15788);
	not 	XG5285 	(g14363,I16521);
	not 	XG5286 	(g12857,I15474);
	not 	XG5287 	(I17989,g14173);
	not 	XG5288 	(I18060,g14198);
	not 	XG5289 	(I18063,g14357);
	not 	XG5290 	(I17956,g14562);
	not 	XG5291 	(I17842,g13051);
	not 	XG5292 	(I17876,g13070);
	not 	XG5293 	(I17916,g13087);
	not 	XG5294 	(I18117,g13302);
	not 	XG5295 	(I17839,g13412);
	not 	XG5296 	(I17754,g13494);
	not 	XG5297 	(g13017,I15633);
	not 	XG5298 	(g13074,I15702);
	not 	XG5299 	(g12977,I15590);
	not 	XG5300 	(g13027,I15647);
	not 	XG5301 	(g13010,I15620);
	not 	XG5302 	(g14252,I16438);
	not 	XG5303 	(g13041,I15667);
	not 	XG5304 	(g13009,I15617);
	not 	XG5305 	(g14330,I16486);
	not 	XG5306 	(g12946,I15564);
	not 	XG5307 	(g13101,I15736);
	not 	XG5308 	(g14383,I16535);
	not 	XG5309 	(g13018,I15636);
	not 	XG5310 	(g14276,I16452);
	not 	XG5311 	(g12978,I15593);
	not 	XG5312 	(g13012,I15626);
	not 	XG5313 	(g13003,I15609);
	not 	XG5314 	(g13055,I15682);
	not 	XG5315 	(g12951,I15569);
	not 	XG5316 	(g13011,I15623);
	not 	XG5317 	(g13075,I15705);
	not 	XG5318 	(g12938,I15556);
	not 	XG5319 	(g13028,I15650);
	not 	XG5320 	(g12918,I15533);
	not 	XG5321 	(g12976,I15587);
	not 	XG5322 	(g11237,I14305);
	not 	XG5323 	(I16489,g12793);
	and 	XG5324 	(g17134,g14851,g5619);
	not 	XG5325 	(g13943,I16231);
	not 	XG5326 	(g10710,I14006);
	not 	XG5327 	(g10851,I14069);
	not 	XG5328 	(g10727,I14016);
	not 	XG5329 	(g10348,I13762);
	not 	XG5330 	(g10347,I13759);
	and 	XG5331 	(g15819,g14101,g3251);
	nand 	XG5332 	(g14107,g11527,g11571);
	nand 	XG5333 	(g14072,g11483,g11571);
	and 	XG5334 	(g16610,g14918,g5260);
	and 	XG5335 	(g15804,g13889,g3223);
	and 	XG5336 	(g14261,g10738,g4507);
	nand 	XG5337 	(g12286,I15130,I15129);
	nand 	XG5338 	(g11761,I14611,I14610);
	not 	XG5339 	(g11705,I14576);
	nor 	XG5340 	(g13603,g10721,g8009);
	not 	XG5341 	(g13574,I16024);
	nand 	XG5342 	(g11906,I14714,I14713);
	nand 	XG5343 	(g12336,I15176,I15175);
	and 	XG5344 	(g16672,g15008,g6295);
	and 	XG5345 	(g17119,g14800,g5272);
	nand 	XG5346 	(g11153,I14206,I14205);
	and 	XG5347 	(g16199,g14051,g3614);
	and 	XG5348 	(g16535,g14848,g5595);
	and 	XG5349 	(g15880,g13980,g3211);
	and 	XG5350 	(g17177,g14984,g6657);
	nor 	XG5351 	(g14320,g11111,g9257);
	and 	XG5352 	(g13853,g10620,g4549);
	nand 	XG5353 	(I17460,g1300,g13378);
	not 	XG5354 	(I15862,g11215);
	nand 	XG5355 	(I15194,I15193,g9935);
	and 	XG5356 	(g15851,g14157,g3953);
	and 	XG5357 	(g12953,g11048,g411);
	and 	XG5358 	(g16705,g15024,g6299);
	nand 	XG5359 	(g11944,I14766,I14765);
	nand 	XG5360 	(g13897,g11519,g3329,g11217,g3211);
	not 	XG5361 	(g11929,I14745);
	and 	XG5362 	(g16593,g14885,g5599);
	and 	XG5363 	(g16673,g14822,g6617);
	nand 	XG5364 	(g17315,g14503,g9516,g9564);
	nor 	XG5365 	(g14522,g12656,g9924);
	nor 	XG5366 	(g14425,g12656,g5644);
	and 	XG5367 	(g15837,g14127,g3255);
	nand 	XG5368 	(g12136,I14993,I14992);
	not 	XG5369 	(g12490,I15316);
	and 	XG5370 	(g15967,g14058,g3913);
	nand 	XG5371 	(g14569,g8481,g3329,g11194,g3195);
	nand 	XG5372 	(g12538,I15335,I15334);
	and 	XG5373 	(g16670,g14999,g5953);
	and 	XG5374 	(g14035,g11048,g699);
	and 	XG5375 	(g15815,g14075,g3594);
	nand 	XG5376 	(g12187,I15043,I15042);
	nor 	XG5377 	(g13004,g10741,g7933);
	nand 	XG5378 	(g11323,I14352,I14351);
	not 	XG5379 	(g13223,I15800);
	or 	XG5380 	(g13969,g8913,g11448);
	nor 	XG5381 	(g14988,g10805,g10812,g10816);
	and 	XG5382 	(g13156,g10805,g10812,g10816);
	not 	XG5383 	(I16593,g10498);
	and 	XG5384 	(g15783,g14098,g3215);
	and 	XG5385 	(g15848,g13892,g3259);
	and 	XG5386 	(g16841,g14858,g5913);
	or 	XG5387 	(g16187,g13486,g8822);
	nor 	XG5388 	(g13539,g12735,g8594);
	and 	XG5389 	(g16516,g14627,g5228);
	not 	XG5390 	(I16163,g11930);
	and 	XG5391 	(g15859,g13923,g3610);
	and 	XG5392 	(g16871,g14908,g6597);
	nor 	XG5393 	(g16424,g13628,g8064);
	and 	XG5394 	(g15793,g13873,g3219);
	and 	XG5395 	(g17057,g13173,g446);
	nand 	XG5396 	(g11559,I14510,I14509);
	and 	XG5397 	(g15818,g14082,g3941);
	not 	XG5398 	(g15568,g14984);
	nand 	XG5399 	(g15030,g12680,g12716);
	not 	XG5400 	(g17791,g14950);
	nand 	XG5401 	(g15011,g12632,g12716);
	nand 	XG5402 	(g15829,g13831,g4112);
	nor 	XG5403 	(g14247,g10869,g9934);
	nand 	XG5404 	(I17446,g956,g13336);
	and 	XG5405 	(g17617,g13326,g7885);
	or 	XG5406 	(I18421,g14395,g14417,g14447);
	nand 	XG5407 	(g13092,g10761,g1061);
	nand 	XG5408 	(g17243,g14212,g7247);
	and 	XG5409 	(g17693,g13291,g1306);
	not 	XG5410 	(g14873,I16898);
	and 	XG5411 	(g16736,g15036,g6303);
	and 	XG5412 	(g16642,g14981,g6633);
	nor 	XG5413 	(g13005,g10762,g7939);
	not 	XG5414 	(I16512,g12811);
	nor 	XG5415 	(g13129,g10762,g7553);
	and 	XG5416 	(g12979,g11048,g424);
	not 	XG5417 	(g13545,I16010);
	and 	XG5418 	(g16532,g14841,g5252);
	and 	XG5419 	(g17784,g13215,g1152);
	and 	XG5420 	(g16596,g14892,g5941);
	not 	XG5421 	(g11720,I14589);
	nand 	XG5422 	(I18680,g14752,g2638);
	not 	XG5423 	(g11845,I14663);
	nand 	XG5424 	(g12431,I15255,I15254);
	or 	XG5425 	(I18492,g14446,g14513,g14538);
	not 	XG5426 	(g14348,g10887);
	not 	XG5427 	(g17777,g14908);
	nand 	XG5428 	(g14978,g10491,g12716);
	not 	XG5429 	(g14785,g12629);
	nand 	XG5430 	(g15045,g7142,g12716);
	nor 	XG5431 	(g14347,g11123,g9309);
	or 	XG5432 	(I18385,g14360,g14391,g14413);
	not 	XG5433 	(g12039,I14899);
	nor 	XG5434 	(g15669,g14272,g11945);
	and 	XG5435 	(g16844,g13000,g7212);
	and 	XG5436 	(g12931,g11048,g392);
	and 	XG5437 	(g15808,g14048,g3590);
	nand 	XG5438 	(I17379,g1129,g13336);
	not 	XG5439 	(g11986,I14830);
	and 	XG5440 	(g16730,g14723,g5212);
	not 	XG5441 	(g11931,I14749);
	nand 	XG5442 	(I14497,g8737,g9020);
	nand 	XG5443 	(g14830,g12721,g6723,g12211,g6605);
	and 	XG5444 	(g13778,g10597,g4540);
	nand 	XG5445 	(g12028,I14885,I14884);
	nor 	XG5446 	(g13377,g10762,g7873);
	and 	XG5447 	(g15823,g14116,g3945);
	not 	XG5448 	(I15869,g11234);
	nor 	XG5449 	(g16292,g13134,g7943);
	nand 	XG5450 	(I15242,I15241,g10003);
	nand 	XG5451 	(g12100,I14957,I14956);
	nand 	XG5452 	(g13968,g11631,g4031,g11255,g3913);
	not 	XG5453 	(I15981,g11290);
	nand 	XG5454 	(g11189,I14249,I14248);
	nand 	XG5455 	(I18633,g14713,g2504);
	not 	XG5456 	(g16305,g13346);
	and 	XG5457 	(g16590,g14683,g5236);
	and 	XG5458 	(g13282,g11480,g3546);
	and 	XG5459 	(g13030,g11048,g429);
	nand 	XG5460 	(g17586,g14601,g14638);
	nand 	XG5461 	(g13139,g10061,g6723,g12137,g6589);
	nor 	XG5462 	(g12980,g10741,g7909);
	not 	XG5463 	(g11855,I14671);
	not 	XG5464 	(g11820,I14644);
	not 	XG5465 	(g11872,I14684);
	not 	XG5466 	(g11894,I14702);
	not 	XG5467 	(g11823,I14647);
	not 	XG5468 	(g11920,I14730);
	not 	XG5469 	(g11897,I14705);
	not 	XG5470 	(g11790,I14630);
	not 	XG5471 	(I16120,g11868);
	nand 	XG5472 	(g11206,I14277,I14276);
	nor 	XG5473 	(g13094,g10762,g7487);
	and 	XG5474 	(g16484,g14755,g5244);
	and 	XG5475 	(g16614,g14933,g5945);
	and 	XG5476 	(g15840,g14142,g3949);
	nand 	XG5477 	(g14946,g12672,g6346,g12173,g6247);
	not 	XG5478 	(g11842,I14660);
	not 	XG5479 	(g10499,I13872);
	and 	XG5480 	(g16483,g14915,g5224);
	not 	XG5481 	(g17718,g14776);
	not 	XG5482 	(g17585,g14974);
	not 	XG5483 	(g17648,g15024);
	not 	XG5484 	(g17505,g14899);
	nor 	XG5485 	(g13044,g10762,g7349);
	not 	XG5486 	(g17521,g14727);
	not 	XG5487 	(g17642,g14691);
	nand 	XG5488 	(g14924,g12505,g12558);
	nand 	XG5489 	(g14882,g12453,g12558);
	not 	XG5490 	(g17498,g14688);
	not 	XG5491 	(g17603,g14993);
	nor 	XG5492 	(g13013,g10762,g7957);
	or 	XG5493 	(g16173,g13464,g8796);
	not 	XG5494 	(g11941,I14761);
	not 	XG5495 	(g11917,I14727);
	not 	XG5496 	(g11875,I14687);
	not 	XG5497 	(g11852,I14668);
	not 	XG5498 	(g14204,g12155);
	or 	XG5499 	(g16926,g11780,g11804,g14061);
	and 	XG5500 	(g16612,g14927,g5603);
	nand 	XG5501 	(g17412,g14489,g14520);
	nor 	XG5502 	(g13325,g10741,g7841);
	nor 	XG5503 	(g13110,g10741,g7841);
	nand 	XG5504 	(g13479,g12526,g12590,g12639,g12686);
	and 	XG5505 	(g16637,g14968,g5949);
	and 	XG5506 	(g13415,g11048,g837);
	nor 	XG5507 	(g13125,g10762,g7863);
	nor 	XG5508 	(g13341,g10762,g7863);
	or 	XG5509 	(g14309,g11048,g10320);
	and 	XG5510 	(g15810,g14055,g3937);
	nor 	XG5511 	(g13114,g10741,g7528);
	not 	XG5512 	(I16596,g12640);
	not 	XG5513 	(g15705,g13217);
	nor 	XG5514 	(g13021,g10741,g7544);
	nand 	XG5515 	(g14014,g11519,g3298,g11217,g3199);
	nand 	XG5516 	(g14422,g8481,g3298,g11194,g3187);
	nand 	XG5517 	(g16757,g11675,g14120,g13886,g13911);
	not 	XG5518 	(g11772,I14623);
	not 	XG5519 	(g11706,I14579);
	or 	XG5520 	(g16876,g11755,g11773,g14028);
	or 	XG5521 	(g16261,g13469,g7898);
	not 	XG5522 	(g11829,I14653);
	not 	XG5523 	(g11900,I14708);
	nor 	XG5524 	(g15647,g14248,g11924);
	not 	XG5525 	(g17741,g12972);
	nand 	XG5526 	(g12436,I15264,I15263);
	not 	XG5527 	(I15834,g11164);
	not 	XG5528 	(g12477,I15295);
	nor 	XG5529 	(g14211,g10823,g9779);
	and 	XG5530 	(g13833,g10613,g4546);
	and 	XG5531 	(g16537,g14855,g5937);
	not 	XG5532 	(g15614,g14914);
	nor 	XG5533 	(g10488,g10336,g7133,g4616);
	not 	XG5534 	(g13414,g11048);
	not 	XG5535 	(g13312,g11048);
	not 	XG5536 	(g14034,g11048);
	not 	XG5537 	(g13305,g11048);
	not 	XG5538 	(g14063,g11048);
	not 	XG5539 	(g14179,g11048);
	not 	XG5540 	(g13458,g11048);
	not 	XG5541 	(g13323,g11048);
	not 	XG5542 	(g13999,g11048);
	not 	XG5543 	(g14032,g11048);
	not 	XG5544 	(g13474,g11048);
	not 	XG5545 	(g14584,g11048);
	not 	XG5546 	(g13334,g11048);
	not 	XG5547 	(g13975,g11048);
	not 	XG5548 	(g14166,g11048);
	not 	XG5549 	(g14065,g11048);
	not 	XG5550 	(I16468,g12760);
	nand 	XG5551 	(g14636,g12563,g5677,g12029,g5595);
	nand 	XG5552 	(g14750,g12721,g6715,g12137,g6633);
	and 	XG5553 	(g16808,g14825,g6653);
	and 	XG5554 	(g17138,g13239,g255);
	nand 	XG5555 	(g12539,I15342,I15341);
	nor 	XG5556 	(g15106,g10430,g12872);
	nor 	XG5557 	(g17213,g13501,g11107);
	and 	XG5558 	(g15872,g14234,g9095);
	nand 	XG5559 	(g11980,I14818,I14817);
	and 	XG5560 	(g16758,g14758,g5220);
	not 	XG5561 	(g14912,I16917);
	not 	XG5562 	(g13267,I15831);
	not 	XG5563 	(g11793,I14633);
	not 	XG5564 	(g11878,I14690);
	not 	XG5565 	(g11826,I14650);
	not 	XG5566 	(g11744,I14602);
	not 	XG5567 	(I16733,g12026);
	and 	XG5568 	(g13737,g10571,g4501);
	not 	XG5569 	(I16538,g10417);
	nand 	XG5570 	(g13104,g10794,g1404);
	and 	XG5571 	(g15912,g14018,g3562);
	and 	XG5572 	(g16185,g14011,g3263);
	not 	XG5573 	(g11317,I14346);
	not 	XG5574 	(g11136,I14192);
	nand 	XG5575 	(g11193,I14259,I14258);
	nor 	XG5576 	(g14437,g11178,g9527);
	or 	XG5577 	(g10589,g7201,g7223);
	and 	XG5578 	(g15995,g10666,g1157,g13314);
	and 	XG5579 	(g15813,g14069,g3247);
	nand 	XG5580 	(I14399,I14398,g8542);
	nand 	XG5581 	(g13907,g11631,g4023,g11225,g3941);
	and 	XG5582 	(g16591,g14879,g5256);
	nand 	XG5583 	(g11511,I14482,I14481);
	and 	XG5584 	(g14216,g10608,g7631);
	not 	XG5585 	(g11966,I14800);
	not 	XG5586 	(g17609,g14817);
	not 	XG5587 	(g17527,g14741);
	not 	XG5588 	(g10363,I13779);
	and 	XG5589 	(g15812,g13915,g3227);
	and 	XG5590 	(g15820,g13955,g3578);
	and 	XG5591 	(g16518,g14956,g5571);
	not 	XG5592 	(I15846,g11183);
	nand 	XG5593 	(g13040,g9780,g5308,g12002,g5196);
	not 	XG5594 	(g10385,I13805);
	or 	XG5595 	(g15727,g11010,g13333,g13345,g13383);
	nand 	XG5596 	(g16663,g12292,g14655,g13834,g13854);
	not 	XG5597 	(I13889,g7598);
	not 	XG5598 	(g11294,g7598);
	nand 	XG5599 	(g17474,g14521,g14547);
	nand 	XG5600 	(I15148,I15147,g9864);
	not 	XG5601 	(g17496,g14683);
	not 	XG5602 	(g17600,g14659);
	nand 	XG5603 	(g14876,g12443,g12492);
	not 	XG5604 	(g18061,g14800);
	nand 	XG5605 	(g14794,g12772,g12492);
	not 	XG5606 	(g17673,g14723);
	not 	XG5607 	(g17414,g14627);
	not 	XG5608 	(g17518,g14918);
	and 	XG5609 	(g13290,g11534,g3897);
	nand 	XG5610 	(g11135,I14187,I14186);
	and 	XG5611 	(g16706,g14868,g6621);
	not 	XG5612 	(g16608,g14116);
	not 	XG5613 	(g16725,g13963);
	not 	XG5614 	(g16529,g14055);
	not 	XG5615 	(g16658,g14157);
	not 	XG5616 	(g17746,g14825);
	not 	XG5617 	(g17721,g12915);
	not 	XG5618 	(g17611,g14822);
	not 	XG5619 	(g17651,g14868);
	nand 	XG5620 	(g13086,g10003,g6346,g12101,g6235);
	not 	XG5621 	(I16492,g12430);
	not 	XG5622 	(g17416,g14956);
	not 	XG5623 	(g17522,g14927);
	nand 	XG5624 	(g14962,g10281,g12558);
	not 	XG5625 	(g17579,g14959);
	nand 	XG5626 	(g14845,g12798,g12558);
	not 	XG5627 	(g17476,g14665);
	nand 	XG5628 	(g12224,I15089,I15088);
	and 	XG5629 	(g14496,I16618,g12197,g12244,g12411);
	nor 	XG5630 	(g13517,g12692,g8541);
	nor 	XG5631 	(g15608,g14212,g11885);
	and 	XG5632 	(g16731,g12941,g7153);
	or 	XG5633 	(I18417,g14392,g14414,g14444);
	and 	XG5634 	(g15861,g14170,g3957);
	not 	XG5635 	(g10384,I13802);
	nand 	XG5636 	(I14369,I14368,g8481);
	nand 	XG5637 	(g13516,g11412,g11444,g11490,g11533);
	nand 	XG5638 	(I14370,I14368,g3303);
	and 	XG5639 	(g13942,g12512,g5897);
	nand 	XG5640 	(g14066,g11473,g11514);
	not 	XG5641 	(g16582,g13915);
	not 	XG5642 	(g16652,g13892);
	not 	XG5643 	(g16522,g13889);
	not 	XG5644 	(g16623,g14127);
	nand 	XG5645 	(g14038,g11435,g11514);
	not 	XG5646 	(g17681,g14735);
	not 	XG5647 	(g17524,g14933);
	not 	XG5648 	(g17479,g14855);
	not 	XG5649 	(g17606,g14999);
	nor 	XG5650 	(g13824,g11702,g8623);
	nor 	XG5651 	(g13772,g11702,g3990);
	not 	XG5652 	(I15811,g11128);
	or 	XG5653 	(I18449,g14415,g14445,g14512);
	not 	XG5654 	(I16471,g12367);
	not 	XG5655 	(g12183,I15033);
	and 	XG5656 	(g17153,g14943,g6311);
	not 	XG5657 	(g13189,g10762);
	not 	XG5658 	(I15821,g11143);
	not 	XG5659 	(g16774,g14024);
	not 	XG5660 	(g17144,g14085);
	and 	XG5661 	(g16704,g15018,g5957);
	or 	XG5662 	(I18452,g14418,g14448,g14514);
	nand 	XG5663 	(I14400,I14398,g3654);
	not 	XG5664 	(g13584,g12735);
	not 	XG5665 	(g13932,g11534);
	not 	XG5666 	(g16773,g14021);
	not 	XG5667 	(g16630,g14142);
	not 	XG5668 	(g16814,g14058);
	not 	XG5669 	(g16589,g14082);
	not 	XG5670 	(g16692,g14170);
	nor 	XG5671 	(g14382,g11139,g9390);
	not 	XG5672 	(g16280,g13330);
	not 	XG5673 	(g15830,g13432);
	not 	XG5674 	(I16676,g10588);
	not 	XG5675 	(I16028,g12381);
	not 	XG5676 	(g14149,g12381);
	not 	XG5677 	(g14205,g12381);
	not 	XG5678 	(I15921,g12381);
	not 	XG5679 	(g14183,g12381);
	not 	XG5680 	(I15954,g12381);
	not 	XG5681 	(g14169,g12381);
	not 	XG5682 	(I15918,g12381);
	not 	XG5683 	(g14150,g12381);
	not 	XG5684 	(I15932,g12381);
	not 	XG5685 	(g14203,g12381);
	not 	XG5686 	(g14191,g12381);
	not 	XG5687 	(g14184,g12381);
	not 	XG5688 	(I15942,g12381);
	not 	XG5689 	(g14219,g12381);
	not 	XG5690 	(g14255,g12381);
	not 	XG5691 	(I15987,g12381);
	nand 	XG5692 	(g12144,I15004,I15003);
	not 	XG5693 	(g13278,g10738);
	not 	XG5694 	(g13061,g10981);
	not 	XG5695 	(g13106,g10981);
	not 	XG5696 	(g13082,g10981);
	not 	XG5697 	(g13484,g10981);
	not 	XG5698 	(g13036,g10981);
	not 	XG5699 	(g13037,g10981);
	not 	XG5700 	(I16610,g10981);
	not 	XG5701 	(g13505,g10981);
	not 	XG5702 	(g13062,g10981);
	not 	XG5703 	(g13522,g10981);
	not 	XG5704 	(I16663,g10981);
	not 	XG5705 	(I15727,g10981);
	not 	XG5706 	(g13117,g10981);
	not 	XG5707 	(I16579,g10981);
	not 	XG5708 	(I16660,g10981);
	not 	XG5709 	(I16688,g10981);
	nand 	XG5710 	(g13498,g12416,g12462,g12522,g12577);
	and 	XG5711 	(g17726,g13315,g1467);
	not 	XG5712 	(I15878,g11249);
	not 	XG5713 	(I16564,g10429);
	not 	XG5714 	(g17612,g15014);
	not 	XG5715 	(g17589,g14981);
	not 	XG5716 	(g15755,g13134);
	not 	XG5717 	(g17473,g14841);
	not 	XG5718 	(g17390,g14755);
	and 	XG5719 	(g16842,g14861,g6279);
	nand 	XG5720 	(g13109,g10003,g6369,g12173,g6279);
	not 	XG5721 	(g17738,g14813);
	not 	XG5722 	(g15479,g14895);
	nand 	XG5723 	(g14803,g12497,g5308,g12059,g5208);
	or 	XG5724 	(g14187,g11771,g8871);
	not 	XG5725 	(g14297,g10869);
	not 	XG5726 	(g17737,g14810);
	not 	XG5727 	(g17583,g14968);
	not 	XG5728 	(g14700,g12512);
	not 	XG5729 	(g17756,g14858);
	not 	XG5730 	(g17645,g15018);
	not 	XG5731 	(g17503,g14892);
	not 	XG5732 	(I16289,g12107);
	not 	XG5733 	(g16030,g13570);
	nand 	XG5734 	(I15166,g9823,g9904);
	nand 	XG5735 	(g14598,g12497,g5331,g12002,g5248);
	not 	XG5736 	(g11987,I14833);
	not 	XG5737 	(g13174,g10741);
	not 	XG5738 	(g15746,g13121);
	and 	XG5739 	(g13974,g12578,g6243);
	and 	XG5740 	(g17771,g13190,g13288);
	not 	XG5741 	(g15756,g13315);
	not 	XG5742 	(g16311,g13273);
	and 	XG5743 	(g15814,g13920,g3574);
	nand 	XG5744 	(I14530,g8873,g8840);
	and 	XG5745 	(g16843,g14864,g6251);
	nand 	XG5746 	(g14088,g11631,g4000,g11255,g3901);
	not 	XG5747 	(I16651,g10542);
	nand 	XG5748 	(I17474,g1105,g13336);
	nor 	XG5749 	(g16581,g8086,g13756);
	not 	XG5750 	(g17735,g14807);
	not 	XG5751 	(g15344,g14851);
	nand 	XG5752 	(g14664,g12497,g5339,g12059,g5220);
	not 	XG5753 	(g16583,g14069);
	nand 	XG5754 	(g14104,g8864,g11514);
	not 	XG5755 	(g16472,g14098);
	not 	XG5756 	(g16509,g13873);
	nand 	XG5757 	(g14005,g11729,g11514);
	not 	XG5758 	(g16602,g14101);
	not 	XG5759 	(I15872,g11236);
	not 	XG5760 	(g16771,g14018);
	not 	XG5761 	(g17124,g14051);
	not 	XG5762 	(g17499,g14885);
	not 	XG5763 	(g17477,g14848);
	not 	XG5764 	(g17762,g13000);
	not 	XG5765 	(g15842,g13469);
	not 	XG5766 	(g16515,g13486);
	not 	XG5767 	(I15814,g11129);
	nand 	XG5768 	(I14211,g9295,g9252);
	not 	XG5769 	(g13555,g12692);
	nand 	XG5770 	(g14136,g8906,g11571);
	not 	XG5771 	(g13901,g11480);
	nand 	XG5772 	(g14045,g11747,g11571);
	not 	XG5773 	(g16743,g13986);
	not 	XG5774 	(g17676,g12941);
	nand 	XG5775 	(I15243,I15241,g6351);
	and 	XG5776 	(g14581,I16695,g12357,g12428,g12587);
	and 	XG5777 	(g16634,g14953,g5264);
	nor 	XG5778 	(g14411,g11160,g9460);
	or 	XG5779 	(g13888,g11691,g2941);
	not 	XG5780 	(I17416,g13806);
	not 	XG5781 	(I15843,g11181);
	not 	XG5782 	(g10473,I13857);
	nand 	XG5783 	(I17883,g1135,g13336);
	nor 	XG5784 	(g14271,g10874,g10002);
	and 	XG5785 	(g15794,g14008,g3239);
	not 	XG5786 	(g12077,I14939);
	nor 	XG5787 	(g12858,g10430,g10365);
	not 	XG5788 	(g12108,I14964);
	not 	XG5789 	(g16689,g13923);
	not 	XG5790 	(g16655,g14151);
	not 	XG5791 	(g16585,g14075);
	not 	XG5792 	(g16527,g14048);
	nand 	XG5793 	(g13515,g12464,g12524,g12588,g12628);
	and 	XG5794 	(g14528,I16646,g12245,g12306,g12459);
	and 	XG5795 	(g14555,I16671,g12307,g12356,g12521);
	not 	XG5796 	(g17759,g14864);
	not 	XG5797 	(g15562,g14943);
	and 	XG5798 	(g13887,g12402,g5204);
	not 	XG5799 	(g15731,g13326);
	nand 	XG5800 	(g17137,g13527,g13511,g13727);
	not 	XG5801 	(g16645,g13756);
	and 	XG5802 	(g16869,g14902,g6259);
	not 	XG5803 	(I15765,g10823);
	not 	XG5804 	(g14238,g10823);
	not 	XG5805 	(g17497,g14879);
	not 	XG5806 	(g14630,g12402);
	not 	XG5807 	(g17389,g14915);
	not 	XG5808 	(g17472,g14656);
	not 	XG5809 	(g17576,g14953);
	not 	XG5810 	(g17707,g14758);
	not 	XG5811 	(I13906,g7620);
	not 	XG5812 	(g11336,g7620);
	not 	XG5813 	(g16482,g13464);
	not 	XG5814 	(g15750,g13291);
	and 	XG5815 	(g16617,g14940,g6287);
	nor 	XG5816 	(g13631,g10733,g8068);
	not 	XG5817 	(g16740,g13980);
	not 	XG5818 	(g17092,g14011);
	nand 	XG5819 	(I15149,I15147,g5659);
	not 	XG5820 	(g16720,g14234);
	not 	XG5821 	(g16523,g14041);
	not 	XG5822 	(g16510,g14008);
	not 	XG5823 	(g16584,g13920);
	not 	XG5824 	(g16605,g13955);
	not 	XG5825 	(g14321,g10874);
	not 	XG5826 	(g17610,g15008);
	not 	XG5827 	(g17758,g14861);
	not 	XG5828 	(g14744,g12578);
	not 	XG5829 	(g17684,g15036);
	not 	XG5830 	(g17774,g14902);
	not 	XG5831 	(g17528,g14940);
	nand 	XG5832 	(g17571,g14367,g8579);
	or 	XG5833 	(g16076,g10736,g13081);
	nand 	XG5834 	(I14428,I14427,g8595);
	nor 	XG5835 	(g17194,g13480,g11039);
	and 	XG5836 	(g15856,g14223,g9056);
	and 	XG5837 	(g15805,g14041,g3243);
	and 	XG5838 	(g16531,g14656,g5232);
	and 	XG5839 	(g15882,g13986,g3554);
	nand 	XG5840 	(g14971,g12581,g12667);
	nand 	XG5841 	(g15027,g10341,g12667);
	nand 	XG5842 	(g13118,g9935,g6031,g12067,g5897);
	nand 	XG5843 	(g14740,g12614,g6031,g12129,g5913);
	and 	XG5844 	(g13321,g11048,g847);
	or 	XG5845 	(g14387,g11048,g9086);
	and 	XG5846 	(g13738,g10572,g8880);
	and 	XG5847 	(g13832,g10612,g8880);
	nand 	XG5848 	(I15195,I15193,g6005);
	nand 	XG5849 	(g12370,I15214,I15213);
	nand 	XG5850 	(g14452,g8542,g3649,g11207,g3538);
	nand 	XG5851 	(g14054,g11576,g3649,g11238,g3550);
	nand 	XG5852 	(I18536,g14642,g2236);
	nor 	XG5853 	(g17420,g14408,g9456);
	nand 	XG5854 	(g12221,I15080,I15079);
	and 	XG5855 	(g16635,g14959,g5607);
	nand 	XG5856 	(g15721,g13385,g311,g7564);
	nand 	XG5857 	(g17312,g14248,g7297);
	nand 	XG5858 	(g13084,g9864,g5677,g12093,g5587);
	and 	XG5859 	(g16759,g14761,g5587);
	nand 	XG5860 	(g14781,g12672,g6377,g12173,g6259);
	nand 	XG5861 	(g13131,g10003,g6377,g12101,g6243);
	and 	XG5862 	(g16702,g14691,g5615);
	and 	XG5863 	(g13633,g10509,g4567);
	nand 	XG5864 	(g14706,g12672,g6369,g12101,g6287);
	and 	XG5865 	(g16047,g10699,g1500,g13322);
	nand 	XG5866 	(g14838,g12405,g12492);
	nand 	XG5867 	(g14921,g10266,g12492);
	and 	XG5868 	(g16519,g14804,g5591);
	and 	XG5869 	(g15821,g14110,g3598);
	nand 	XG5870 	(g14517,g8481,g3321,g11217,g3231);
	nand 	XG5871 	(g13866,g11519,g3321,g11194,g3239);
	nand 	XG5872 	(g16282,g12088,g13939,g4933);
	and 	XG5873 	(g16639,g14974,g6291);
	and 	XG5874 	(g16760,g14764,g5559);
	and 	XG5875 	(g17418,g14407,g9618);
	and 	XG5876 	(g17682,g14637,g9742);
	and 	XG5877 	(g16245,g14708,g14278);
	nand 	XG5878 	(g17748,g12323,g14708,g562);
	and 	XG5879 	(g16804,g14813,g5905);
	nor 	XG5880 	(g13335,g10741,g7851);
	and 	XG5881 	(g17753,g13175,g13281);
	nor 	XG5882 	(g16066,g13307,g10929);
	nor 	XG5883 	(g15992,g13846,g10929);
	nor 	XG5884 	(g16027,g13260,g10929);
	and 	XG5885 	(g15786,g11233,g13940);
	and 	XG5886 	(g16190,g11810,g14626);
	nand 	XG5887 	(g13097,g9780,g5339,g12002,g5204);
	and 	XG5888 	(g15850,g14151,g3606);
	and 	XG5889 	(g15796,g14015,g3586);
	and 	XG5890 	(g16176,g11779,g14596);
	and 	XG5891 	(g15779,g11214,g13909);
	and 	XG5892 	(g15807,g13898,g3570);
	nand 	XG5893 	(g15591,g13202,g4322,g4332);
	nor 	XG5894 	(g14529,g12749,g6336);
	nor 	XG5895 	(g14575,g12749,g10050);
	and 	XG5896 	(g16805,g12972,g7187);
	nor 	XG5897 	(g13622,g11166,g278);
	and 	XG5898 	(g13697,g8608,g11166);
	and 	XG5899 	(g16233,g14251,g6137);
	or 	XG5900 	(g16866,g11044,g13492);
	nand 	XG5901 	(I15106,I15105,g9780);
	and 	XG5902 	(g17405,g13137,g1422);
	and 	XG5903 	(g17321,g13105,g1418);
	and 	XG5904 	(g16513,g13708,g8345);
	nor 	XG5905 	(g13031,g10741,g7301);
	nand 	XG5906 	(g14854,g12563,g5654,g12093,g5555);
	and 	XG5907 	(g13319,g8757,g10658,g8812,g4076);
	and 	XG5908 	(g17469,g13217,g4076);
	nor 	XG5909 	(g15825,g13217,g7666);
	or 	XG5910 	(g16811,g13914,g8690);
	and 	XG5911 	(g15914,g14024,g3905);
	nand 	XG5912 	(g16728,g11639,g14089,g13870,g13884);
	nand 	XG5913 	(g13100,g10061,g6692,g12137,g6581);
	nand 	XG5914 	(g14987,g12721,g6692,g12211,g6593);
	nand 	XG5915 	(I15107,I15105,g5313);
	and 	XG5916 	(g16422,g13627,g8216);
	and 	XG5917 	(g17810,g13246,g1495);
	and 	XG5918 	(g17719,g14675,g9818);
	or 	XG5919 	(g15803,g10528,g12924);
	nand 	XG5920 	(g14696,g12563,g5685,g12093,g5567);
	and 	XG5921 	(g16802,g14807,g5567);
	and 	XG5922 	(g16616,g14741,g6267);
	and 	XG5923 	(g15704,g13504,g3440);
	nor 	XG5924 	(g16090,g13315,g10961);
	nor 	XG5925 	(g16072,g13273,g10961);
	and 	XG5926 	(g17146,g14895,g5965);
	or 	XG5927 	(g15792,g10501,g12920);
	nor 	XG5928 	(g15594,g7285,g13026,g10614);
	nand 	XG5929 	(g13098,g9935,g6023,g12129,g5933);
	and 	XG5930 	(g16803,g14810,g5933);
	and 	XG5931 	(g15749,g13273,g1454);
	or 	XG5932 	(g16970,g11163,g13567);
	nand 	XG5933 	(I15288,I15287,g10061);
	not 	XG5934 	(g16512,g14015);
	not 	XG5935 	(g16626,g14133);
	not 	XG5936 	(g16526,g13898);
	not 	XG5937 	(g16742,g13983);
	not 	XG5938 	(g16606,g14110);
	not 	XG5939 	(g16511,g14130);
	nand 	XG5940 	(g16281,g12054,g13937,g4754);
	and 	XG5941 	(g15841,g13868,g4273);
	nand 	XG5942 	(g12066,I14925,I14924);
	or 	XG5943 	(g16258,g10856,g13247);
	nand 	XG5944 	(g16296,g13501,g9360);
	and 	XG5945 	(g16669,g14993,g5611);
	nand 	XG5946 	(g13499,g11382,g11410,g11442,g11479);
	and 	XG5947 	(g15784,g13977,g3235);
	and 	XG5948 	(g13808,g10607,g4543);
	nand 	XG5949 	(g12191,I15053,I15052);
	nand 	XG5950 	(g17596,g14367,g8686);
	nor 	XG5951 	(g16288,g417,g13794);
	nand 	XG5952 	(g14123,g10928,g10685);
	and 	XG5953 	(g13320,g11048,g417);
	and 	XG5954 	(g10543,g437,g8238);
	and 	XG5955 	(g13299,g11048,g437);
	nand 	XG5956 	(g14898,g12614,g6000,g12129,g5901);
	and 	XG5957 	(g16208,g14085,g3965);
	nand 	XG5958 	(g14570,g8595,g4023,g11255,g3933);
	and 	XG5959 	(g15913,g14021,g3933);
	not 	XG5960 	(g16684,g14223);
	nor 	XG5961 	(g16268,g13121,g7913);
	and 	XG5962 	(g16243,g14275,g6483);
	nand 	XG5963 	(g13069,g9935,g6000,g12067,g5889);
	and 	XG5964 	(g13604,g10487,g4495);
	not 	XG5965 	(g16473,g13977);
	not 	XG5966 	(g16717,g13951);
	not 	XG5967 	(g16716,g13948);
	not 	XG5968 	(g13876,g11432);
	not 	XG5969 	(g13530,g12641);
	nand 	XG5970 	(g11224,I14291,I14290);
	nand 	XG5971 	(g14674,g12614,g6023,g12067,g5941);
	nor 	XG5972 	(g13076,g10741,g7443);
	nand 	XG5973 	(g17364,g14367,g8639);
	nand 	XG5974 	(g14590,g8542,g3680,g11207,g3546);
	nand 	XG5975 	(g13928,g11576,g3680,g11238,g3562);
	and 	XG5976 	(g16674,g15014,g6637);
	and 	XG5977 	(g17401,g13143,g1083);
	and 	XG5978 	(g16764,g14776,g6307);
	nand 	XG5979 	(g17493,g14367,g8659);
	nor 	XG5980 	(g13056,g10741,g7400);
	and 	XG5981 	(g13830,I16143,g11395,g11424,g11543);
	nand 	XG5982 	(g13108,g9864,g5685,g12029,g5551);
	and 	XG5983 	(g13912,g12450,g5551);
	nand 	XG5984 	(g16260,g12088,g13910,g4888);
	nand 	XG5985 	(g16696,g12340,g14682,g13855,g13871);
	or 	XG5986 	(g15732,g11016,g13349,g13384,g13411);
	nand 	XG5987 	(g17363,g14367,g8635);
	and 	XG5988 	(g13042,g11048,g433);
	and 	XG5989 	(g17655,g13342,g7897);
	not 	XG5990 	(g15740,g13342);
	nand 	XG5991 	(g13050,g9864,g5654,g12029,g5543);
	and 	XG5992 	(g16734,g14735,g5961);
	nand 	XG5993 	(g14519,g8595,g4000,g11225,g3889);
	and 	XG5994 	(g16619,g14947,g6629);
	and 	XG5995 	(g16986,g13142,g246);
	nand 	XG5996 	(g13529,g11446,g11492,g11544,g11590);
	and 	XG5997 	(g13671,g10532,g4498);
	nor 	XG5998 	(g13661,g11185,g528);
	nor 	XG5999 	(g13698,g11185,g12527,g528);
	nand 	XG6000 	(g13067,g9780,g5331,g12059,g5240);
	and 	XG6001 	(g16930,g13132,g239);
	and 	XG6002 	(g17643,g14599,g9681);
	nand 	XG6003 	(g13882,g11576,g3672,g11207,g3590);
	nand 	XG6004 	(g14542,g8542,g3672,g11238,g3582);
	and 	XG6005 	(g17424,g13176,g1426);
	or 	XG6006 	(g16506,g10966,g13294);
	and 	XG6007 	(g17480,g14433,g9683);
	and 	XG6008 	(g16766,g12915,g6649);
	nand 	XG6009 	(I14330,g9966,g225);
	and 	XG6010 	(g17123,g13209,g225);
	and 	XG6011 	(g13807,g10606,g4504);
	nand 	XG6012 	(g14930,g12515,g12609);
	nand 	XG6013 	(g15002,g10312,g12609);
	nor 	XG6014 	(g17284,g14317,g9253);
	and 	XG6015 	(g16592,g14688,g5579);
	nor 	XG6016 	(g15628,g14228,g11907);
	and 	XG6017 	(g16761,g12947,g7170);
	not 	XG6018 	(g17713,g12947);
	and 	XG6019 	(g16536,g14996,g5917);
	nand 	XG6020 	(g11962,I14790,I14789);
	nand 	XG6021 	(I14429,I14427,g4005);
	nand 	XG6022 	(I17494,g1448,g13378);
	nand 	XG6023 	(I18587,g14679,g2370);
	not 	XG6024 	(g17672,g14720);
	not 	XG6025 	(g17415,g14797);
	or 	XG6026 	(g16239,g13432,g7892);
	and 	XG6027 	(g15875,g13963,g3961);
	and 	XG6028 	(g17654,g13284,g962);
	nand 	XG6029 	(g13119,g10061,g6715,g12211,g6625);
	and 	XG6030 	(g16870,g14905,g6625);
	nor 	XG6031 	(g14497,g12705,g5990);
	nor 	XG6032 	(g14549,g12705,g9992);
	nor 	XG6033 	(g13078,g10762,g7446);
	nor 	XG6034 	(g15585,g14194,g11862);
	and 	XG6035 	(g16699,g12933,g7134);
	or 	XG6036 	(g15965,g10675,g13035);
	or 	XG6037 	(g16867,g11045,g13493);
	nor 	XG6038 	(g13700,g11615,g3288);
	nor 	XG6039 	(g13765,g11615,g8531);
	nor 	XG6040 	(g14399,g12598,g5297);
	nand 	XG6041 	(g13462,g12294,g12342,g12412,g12449);
	nor 	XG6042 	(g14490,g12598,g9853);
	and 	XG6043 	(g16690,g13867,g8399);
	nor 	XG6044 	(g13032,g10762,g7577);
	and 	XG6045 	(g17307,g14343,g9498);
	and 	XG6046 	(g16221,g14231,g5791);
	and 	XG6047 	(g16737,g15042,g6645);
	nand 	XG6048 	(g14113,g11537,g11626);
	nand 	XG6049 	(g14160,g8958,g11626);
	nor 	XG6050 	(g17239,g13518,g11119);
	and 	XG6051 	(g15883,g14258,g9180);
	and 	XG6052 	(g16534,g14665,g5575);
	not 	XG6053 	(g16746,g14258);
	and 	XG6054 	(g15809,g14154,g3917);
	nand 	XG6055 	(g12969,g10476,g7178,g4388);
	and 	XG6056 	(g16671,g14817,g6275);
	nand 	XG6057 	(g13066,g10590,g7178,g4430);
	and 	XG6058 	(g16653,g13850,g8343);
	and 	XG6059 	(g17149,g13255,g232);
	and 	XG6060 	(g16667,g14659,g5268);
	and 	XG6061 	(g17601,g14572,g9616);
	and 	XG6062 	(g13313,g11048,g475);
	nand 	XG6063 	(g14889,g12824,g12609);
	nand 	XG6064 	(g14965,g12571,g12609);
	or 	XG6065 	(g16022,g10707,g13048);
	and 	XG6066 	(g13771,I16111,g11302,g11355,g11441);
	nor 	XG6067 	(g13730,g11663,g3639);
	nor 	XG6068 	(g13799,g11663,g8584);
	or 	XG6069 	(g16021,g10706,g13047);
	and 	XG6070 	(g15712,g13521,g3791);
	and 	XG6071 	(g16965,g13140,g269);
	and 	XG6072 	(g13020,g11048,g401);
	and 	XG6073 	(g13306,g11048,g441);
	and 	XG6074 	(g17574,g14546,g9554);
	and 	XG6075 	(g16211,g14215,g5445);
	nand 	XG6076 	(g11561,I14518,I14517);
	not 	XG6077 	(g17417,g14804);
	not 	XG6078 	(g17710,g14764);
	not 	XG6079 	(g17709,g14761);
	not 	XG6080 	(g14668,g12450);
	not 	XG6081 	(g14262,g10838);
	and 	XG6082 	(g17769,g13188,g1146);
	nand 	XG6083 	(g14079,g11763,g11626);
	nand 	XG6084 	(g14139,g11584,g11626);
	nor 	XG6085 	(g16313,g13600,g8005);
	nand 	XG6086 	(I17404,g1472,g13378);
	or 	XG6087 	(g14583,g542,g10685);
	or 	XG6088 	(g16882,g11114,g13508);
	not 	XG6089 	(g16290,g13260);
	not 	XG6090 	(g16182,g13846);
	not 	XG6091 	(g15747,g13307);
	and 	XG6092 	(g12939,g11048,g405);
	and 	XG6093 	(g17506,g14505,g9744);
	nand 	XG6094 	(g17246,g14405,g9379,g9439);
	nand 	XG6095 	(g16259,g12054,g13908,g4743);
	and 	XG6096 	(g13029,g11030,g8359);
	or 	XG6097 	(g11737,g8292,g8359);
	and 	XG6098 	(g16707,g15033,g6641);
	and 	XG6099 	(g13564,g12820,g4480);
	and 	XG6100 	(g17391,g14378,g9556);
	and 	XG6101 	(g16638,g14773,g6271);
	nand 	XG6102 	(g17500,g14548,g14573);
	and 	XG6103 	(g17317,g13124,g1079);
	and 	XG6104 	(g17292,g13093,g1075);
	nor 	XG6105 	(g14306,g10887,g10060);
	and 	XG6106 	(g16896,g13120,g262);
	nand 	XG6107 	(g15005,g12622,g12667);
	nand 	XG6108 	(g14937,g10421,g12667);
	not 	XG6109 	(g17504,g15021);
	not 	XG6110 	(g17584,g14773);
	not 	XG6111 	(g17189,g14708);
	or 	XG6112 	(g16052,g10724,g13060);
	nor 	XG6113 	(g17309,g14344,g9305);
	and 	XG6114 	(g13393,g11048,g703);
	nand 	XG6115 	(g10472,I13852,I13851);
	not 	XG6116 	(g15739,g13284);
	nand 	XG6117 	(g16306,g12088,g13971,g4944);
	or 	XG6118 	(g16839,g11035,g13473);
	nand 	XG6119 	(g13083,g4434,g10590,g4392);
	nand 	XG6120 	(g11169,I14230,I14229);
	nand 	XG6121 	(g16586,g13823,g13851);
	or 	XG6122 	(g13526,g301,g10685,g209);
	nor 	XG6123 	(g15754,g13385,g7440,g341);
	not 	XG6124 	(g17523,g14732);
	not 	XG6125 	(g17478,g14996);
	not 	XG6126 	(g17582,g14768);
	not 	XG6127 	(g17502,g14697);
	and 	XG6128 	(g16641,g14782,g6613);
	and 	XG6129 	(g13497,g12155,g2724);
	nor 	XG6130 	(g14291,g12155,g9839);
	nand 	XG6131 	(g15715,g13385,g305,g336);
	not 	XG6132 	(g15831,g13385);
	nand 	XG6133 	(I18579,g14678,g1945);
	nand 	XG6134 	(I17923,g1478,g13378);
	not 	XG6135 	(g16528,g14154);
	not 	XG6136 	(g16588,g13929);
	not 	XG6137 	(g16607,g13960);
	not 	XG6138 	(g16629,g13990);
	not 	XG6139 	(g14639,I16747);
	not 	XG6140 	(g13437,I15937);
	nand 	XG6141 	(g16524,g13798,g13822);
	nand 	XG6142 	(g16299,g13706,g8112,g8160);
	nand 	XG6143 	(I15289,I15287,g6697);
	and 	XG6144 	(g16303,g12921,g4527);
	nand 	XG6145 	(g16507,g13764,g13797);
	nor 	XG6146 	(g17482,g14434,g9523);
	not 	XG6147 	(g15655,g13202);
	not 	XG6148 	(g17811,g12925);
	and 	XG6149 	(g15707,g13506,g4082);
	nand 	XG6150 	(g11923,I14735,I14734);
	nor 	XG6151 	(g14556,g12790,g6682);
	nor 	XG6152 	(g14602,g12790,g10099);
	nand 	XG6153 	(g17220,g14376,g9298,g9369);
	nand 	XG6154 	(g12285,I15123,I15122);
	or 	XG6155 	(I18543,g14516,g14540,g14568);
	and 	XG6156 	(g13461,g11819,g2719);
	and 	XG6157 	(g16611,g14727,g5583);
	and 	XG6158 	(g16598,g14899,g6283);
	nand 	XG6159 	(g17396,g14272,g7345);
	nand 	XG6160 	(g16321,g12088,g13996,g4955);
	not 	XG6161 	(g13249,g10590);
	not 	XG6162 	(g13222,g10590);
	nand 	XG6163 	(g17492,g14367,g8655);
	nand 	XG6164 	(g12592,I15365,I15364);
	or 	XG6165 	(g13858,g10685,g209);
	and 	XG6166 	(g16618,g15039,g6609);
	or 	XG6167 	(I18495,g14449,g14515,g14539);
	and 	XG6168 	(g13998,g12629,g6589);
	nand 	XG6169 	(g17399,g14535,g9574,g9626);
	or 	XG6170 	(g16883,g11115,g13509);
	nand 	XG6171 	(g12999,g4401,g10476,g4392);
	and 	XG6172 	(g14681,g10476,g4392);
	and 	XG6173 	(g14719,g10830,g4392);
	and 	XG6174 	(g14654,g10476,g7178);
	not 	XG6175 	(g13463,g10476);
	not 	XG6176 	(g13107,g10476);
	not 	XG6177 	(g13485,g10476);
	not 	XG6178 	(g13065,g10476);
	or 	XG6179 	(g16959,g11142,g13542);
	not 	XG6180 	(I16755,g12377);
	not 	XG6181 	(g14714,g11405);
	not 	XG6182 	(g14541,g11405);
	not 	XG6183 	(g14833,g11405);
	and 	XG6184 	(g16885,g14950,g6605);
	nand 	XG6185 	(g12482,I15308,I15307);
	or 	XG6186 	(g16448,g10934,g13287);
	not 	XG6187 	(g17637,g12933);
	not 	XG6188 	(g17529,g15039);
	not 	XG6189 	(g17776,g14905);
	not 	XG6190 	(g17652,g15033);
	not 	XG6191 	(g17588,g14782);
	not 	XG6192 	(g17530,g14947);
	not 	XG6193 	(g17687,g15042);
	nand 	XG6194 	(I18485,g14611,g1677);
	and 	XG6195 	(g15700,g13483,g3089);
	and 	XG6196 	(g16202,g14197,g86);
	nand 	XG6197 	(g17595,g14367,g8616);
	or 	XG6198 	(g15910,g10654,g13025);
	nand 	XG6199 	(g13478,g12344,g12414,g12460,g12511);
	or 	XG6200 	(g16928,g11127,g13525);
	nand 	XG6201 	(g12478,I15300,I15299);
	and 	XG6202 	(g14608,I16721,g12429,g12476,g12638);
	nand 	XG6203 	(g12001,I14855,I14854);
	or 	XG6204 	(g16800,g11027,g13436);
	and 	XG6205 	(g13221,g11425,g6946);
	or 	XG6206 	(g14511,g546,g10685);
	nand 	XG6207 	(g17525,g14574,g14600);
	nand 	XG6208 	(g17225,g14367,g8612);
	not 	XG6209 	(g16075,g13597);
	or 	XG6210 	(g16927,g11126,g13524);
	nand 	XG6211 	(g11118,I14171,I14170);
	or 	XG6212 	(g15968,g10677,g13038);
	not 	XG6213 	(g17494,g14339);
	not 	XG6214 	(g17467,g14339);
	or 	XG6215 	(g14977,g8703,g10776);
	or 	XG6216 	(g14078,g8703,g10776);
	or 	XG6217 	(g15017,g8703,g10776);
	or 	XG6218 	(g14936,g8703,g10776);
	or 	XG6219 	(g14888,g8703,g10776);
	or 	XG6220 	(g14044,g8703,g10776);
	or 	XG6221 	(g14844,g8703,g10776);
	or 	XG6222 	(g14119,g8703,g10776);
	not 	XG6223 	(g17573,g12911);
	and 	XG6224 	(g15678,g13846,g1094);
	and 	XG6225 	(g15574,g13202,g4311);
	nand 	XG6226 	(g15710,g13385,g319);
	nand 	XG6227 	(g16278,g13664,g8057,g8102);
	nand 	XG6228 	(g16238,g12054,g13883,g4698);
	nand 	XG6229 	(I18625,g14712,g2079);
	nor 	XG6230 	(g16476,g13667,g8119);
	and 	XG6231 	(g15738,g13260,g1111);
	and 	XG6232 	(g13277,g11432,g3195);
	nor 	XG6233 	(g17198,g14279,g9282);
	nor 	XG6234 	(g17190,g14279,g723);
	nor 	XG6235 	(g17393,g14379,g9386);
	and 	XG6236 	(g16517,g14797,g5248);
	nand 	XG6237 	(g17217,g14194,g7239);
	or 	XG6238 	(g15582,g12925,g8977);
	nand 	XG6239 	(I18529,g14640,g1811);
	and 	XG6240 	(g15817,g13929,g3921);
	and 	XG6241 	(g16595,g14697,g5921);
	and 	XG6242 	(g16324,g182,g13657);
	or 	XG6243 	(g16430,g13657,g182);
	and 	XG6244 	(g16597,g15021,g6263);
	nand 	XG6245 	(g16304,g12054,g13970,g4765);
	and 	XG6246 	(g15822,g13960,g3925);
	and 	XG6247 	(g14193,g10590,g7178);
	and 	XG6248 	(g14210,g10590,g4392);
	and 	XG6249 	(g17692,g13307,g1124);
	and 	XG6250 	(g16613,g14732,g5925);
	nor 	XG6251 	(g14227,g10838,g9863);
	and 	XG6252 	(g15839,g13990,g3929);
	nor 	XG6253 	(g15508,g14279,g10320);
	nor 	XG6254 	(g15372,g14279,g817);
	and 	XG6255 	(g16636,g14768,g5929);
	nor 	XG6256 	(g13500,g12641,g8480);
	and 	XG6257 	(g17786,g13216,g1489);
	and 	XG6258 	(g16621,g13821,g8278);
	and 	XG6259 	(g16474,g13666,g8280);
	and 	XG6260 	(g16729,g14720,g5240);
	and 	XG6261 	(g17156,g13385,g305);
	nand 	XG6262 	(g16316,g13518,g9429);
	nand 	XG6263 	(g16275,g13480,g9291);
	nor 	XG6264 	(g17174,g14279,g9194);
	nor 	XG6265 	(g17148,g14279,g827);
	nand 	XG6266 	(g16319,g13736,g8170,g8224);
	nand 	XG6267 	(g17287,g14228,g7262);
	and 	XG6268 	(g15871,g13951,g3203);
	nand 	XG6269 	(g17290,g14431,g9449,g9506);
	and 	XG6270 	(g15881,g13983,g3582);
	and 	XG6271 	(g15838,g14133,g3602);
	nand 	XG6272 	(g14625,g8595,g4031,g11225,g3897);
	nor 	XG6273 	(g13670,g10756,g8123);
	nor 	XG6274 	(g15170,g14279,g7118);
	nor 	XG6275 	(g17954,g14279,g832);
	and 	XG6276 	(g13805,I16129,g11356,g11394,g11489);
	and 	XG6277 	(g15870,g13948,g3231);
	nor 	XG6278 	(g16044,g13861,g10961);
	not 	XG6279 	(g16197,g13861);
	nor 	XG6280 	(g15578,g14279,g7216);
	nor 	XG6281 	(g15570,g14279,g822);
	and 	XG6282 	(g15795,g14130,g3566);
	and 	XG6283 	(g13656,g11144,g278);
	and 	XG6284 	(g15699,g13861,g1437);
	and 	XG6285 	(g15117,g14454,g4300);
	nor 	XG6286 	(g15120,g13605,g12873);
	nor 	XG6287 	(g15123,g13605,g6975);
	nor 	XG6288 	(g15122,g13605,g6959);
	and 	XG6289 	(g15103,g14454,g4180);
	and 	XG6290 	(g15114,g14454,g4239);
	and 	XG6291 	(g15112,g14454,g4284);
	nor 	XG6292 	(g15061,g13394,g6815);
	and 	XG6293 	(g15118,g14454,g4253);
	nor 	XG6294 	(g15069,g13416,g6828);
	and 	XG6295 	(g15083,g12983,g10362);
	nor 	XG6296 	(g15131,g13638,g12881);
	nor 	XG6297 	(g15146,g7003,g13716);
	nor 	XG6298 	(g15149,g12894,g13745);
	and 	XG6299 	(g15082,g12983,g2697);
	nor 	XG6300 	(g15098,g6927,g13191);
	nor 	XG6301 	(g15057,g13350,g6810);
	and 	XG6302 	(g15075,g12955,g12850);
	nor 	XG6303 	(g15150,g13745,g12895);
	nor 	XG6304 	(g15156,g7050,g13782);
	and 	XG6305 	(g15107,g14454,g4258);
	nor 	XG6306 	(g15143,g13680,g6998);
	nor 	XG6307 	(g17657,g12955,g14751);
	nor 	XG6308 	(g15065,g12840,g13394);
	and 	XG6309 	(g15080,g12983,g12855);
	nor 	XG6310 	(g15062,g13394,g6817);
	nor 	XG6311 	(g15138,g6993,g13680);
	nor 	XG6312 	(g15051,g13350,g6801);
	nor 	XG6313 	(g15070,g13416,g6829);
	nor 	XG6314 	(g15147,g12892,g13716);
	nor 	XG6315 	(g15089,g12861,g13144);
	and 	XG6316 	(g15081,g12983,g2689);
	nor 	XG6317 	(g15068,g13416,g6826);
	and 	XG6318 	(g15113,g14454,g4291);
	and 	XG6319 	(g15110,g14454,g4245);
	nor 	XG6320 	(g17727,g12983,g12486);
	nor 	XG6321 	(g15054,g13350,g12837);
	nor 	XG6322 	(g17694,g12955,g12435);
	nor 	XG6323 	(g15148,g12893,g13716);
	nor 	XG6324 	(g15073,g13416,g12844);
	and 	XG6325 	(g15119,g14454,g4249);
	and 	XG6326 	(g15077,g12955,g2138);
	nor 	XG6327 	(g15128,g12880,g13638);
	nor 	XG6328 	(g15050,g13350,g12834);
	nor 	XG6329 	(g15137,g13680,g6992);
	nor 	XG6330 	(g15164,g12906,g13835);
	and 	XG6331 	(g15115,g14454,g2946);
	nor 	XG6332 	(g15097,g13191,g12868);
	nor 	XG6333 	(g15129,g13638,g6984);
	nor 	XG6334 	(g15121,g13605,g12874);
	and 	XG6335 	(g18655,g14454,g15106);
	nor 	XG6336 	(g15067,g13394,g12842);
	nor 	XG6337 	(g15074,g13416,g12845);
	or 	XG6338 	(g15124,g4581,g13605);
	nor 	XG6339 	(g15049,g6799,g13350);
	nor 	XG6340 	(g15165,g13835,g12907);
	nor 	XG6341 	(g15056,g13350,g6809);
	nor 	XG6342 	(g15066,g13394,g12841);
	nor 	XG6343 	(g15087,g13144,g12860);
	nor 	XG6344 	(g15141,g13680,g12888);
	and 	XG6345 	(g15079,g12955,g2151);
	nor 	XG6346 	(g15100,g12870,g13191);
	or 	XG6347 	(g15125,g13605,g10363);
	nor 	XG6348 	(g15053,g13350,g12836);
	nor 	XG6349 	(g15071,g13416,g6831);
	and 	XG6350 	(g15084,g12983,g2710);
	nor 	XG6351 	(g15132,g13638,g12882);
	nor 	XG6352 	(g15126,g13605,g12878);
	nor 	XG6353 	(g15130,g6985,g13638);
	nor 	XG6354 	(g17619,g12955,g10179);
	nor 	XG6355 	(g15152,g12896,g13745);
	nor 	XG6356 	(g15099,g12869,g13191);
	nor 	XG6357 	(g15091,g12863,g13177);
	nor 	XG6358 	(g15092,g13177,g12864);
	nor 	XG6359 	(g15096,g12867,g13191);
	and 	XG6360 	(g15076,g12955,g2130);
	nor 	XG6361 	(g17700,g12983,g14792);
	nor 	XG6362 	(g15090,g12862,g13144);
	nor 	XG6363 	(g15160,g13809,g12903);
	nor 	XG6364 	(g15157,g12900,g13782);
	nor 	XG6365 	(g15144,g12890,g13716);
	and 	XG6366 	(g15078,g12955,g10361);
	nor 	XG6367 	(g15086,g12859,g13144);
	nor 	XG6368 	(g15142,g12889,g13680);
	nor 	XG6369 	(g15154,g12898,g13782);
	nor 	XG6370 	(g15134,g12884,g13638);
	nor 	XG6371 	(g15127,g13605,g12879);
	nor 	XG6372 	(g15060,g6814,g13350);
	nor 	XG6373 	(g15166,g7096,g13835);
	nor 	XG6374 	(g15102,g6954,g14591);
	and 	XG6375 	(g15116,g14454,g4297);
	and 	XG6376 	(g15111,g14454,g4281);
	nor 	XG6377 	(g15139,g13680,g12886);
	nor 	XG6378 	(g15151,g7027,g13745);
	nor 	XG6379 	(g15161,g7073,g13809);
	nor 	XG6380 	(g15064,g13394,g6820);
	nor 	XG6381 	(g15167,g12908,g13835);
	nor 	XG6382 	(g15155,g13782,g12899);
	nor 	XG6383 	(g15093,g6904,g13177);
	nor 	XG6384 	(g15088,g6874,g13144);
	and 	XG6385 	(g15109,g14454,g4269);
	nor 	XG6386 	(g15072,g12843,g13416);
	and 	XG6387 	(g15104,g14454,g6955);
	nor 	XG6388 	(g15133,g13638,g12883);
	nor 	XG6389 	(g15135,g13638,g6990);
	nor 	XG6390 	(g15095,g12866,g13177);
	nor 	XG6391 	(g15153,g12897,g13745);
	nor 	XG6392 	(g15094,g12865,g13177);
	nor 	XG6393 	(g15101,g14591,g12871);
	nor 	XG6394 	(g15058,g13350,g12838);
	nor 	XG6395 	(g15055,g13350,g6808);
	nor 	XG6396 	(g15162,g12904,g13809);
	nor 	XG6397 	(g15145,g13716,g12891);
	nor 	XG6398 	(g15159,g12902,g13809);
	nor 	XG6399 	(g15059,g13350,g12839);
	nor 	XG6400 	(g15158,g12901,g13782);
	nor 	XG6401 	(g15140,g13680,g12887);
	nor 	XG6402 	(g15163,g12905,g13809);
	and 	XG6403 	(g15108,g14454,g4264);
	nor 	XG6404 	(g15168,g12909,g13835);
	nor 	XG6405 	(g15052,g13350,g12835);
	nor 	XG6406 	(g17663,g12983,g10205);
	and 	XG6407 	(g15105,g14454,g4235);
	nor 	XG6408 	(g15136,g12885,g13680);
	nor 	XG6409 	(g15063,g13394,g6818);
	not 	XG6410 	(I18301,g12976);
	not 	XG6411 	(I18214,g12918);
	not 	XG6412 	(I18446,g13028);
	not 	XG6413 	(I18248,g12938);
	not 	XG6414 	(I18574,g13075);
	not 	XG6415 	(I18373,g13011);
	not 	XG6416 	(I18280,g12951);
	not 	XG6417 	(I18526,g13055);
	not 	XG6418 	(I18344,g13003);
	not 	XG6419 	(I18379,g13012);
	not 	XG6420 	(I18310,g12978);
	not 	XG6421 	(I17653,g14276);
	not 	XG6422 	(I18411,g13018);
	not 	XG6423 	(I17750,g14383);
	not 	XG6424 	(I18674,g13101);
	not 	XG6425 	(I18259,g12946);
	not 	XG6426 	(I17695,g14330);
	not 	XG6427 	(I18364,g13009);
	not 	XG6428 	(I18479,g13041);
	not 	XG6429 	(I17636,g14252);
	not 	XG6430 	(I18367,g13010);
	not 	XG6431 	(I18443,g13027);
	not 	XG6432 	(I18307,g12977);
	not 	XG6433 	(I18571,g13074);
	not 	XG6434 	(I18408,g13017);
	not 	XG6435 	(g16580,I17754);
	not 	XG6436 	(g16643,I17839);
	not 	XG6437 	(g16963,I18117);
	not 	XG6438 	(g16708,I17916);
	not 	XG6439 	(g16676,I17876);
	not 	XG6440 	(g16644,I17842);
	not 	XG6441 	(g16738,I17956);
	not 	XG6442 	(g16873,I18063);
	not 	XG6443 	(g16872,I18060);
	not 	XG6444 	(g16767,I17989);
	not 	XG6445 	(I17008,g12857);
	not 	XG6446 	(I17118,g14363);
	not 	XG6447 	(I18168,g13191);
	not 	XG6448 	(I18177,g13191);
	not 	XG6449 	(I18270,g13191);
	not 	XG6450 	(I18125,g13191);
	not 	XG6451 	(I17763,g13191);
	not 	XG6452 	(g17471,g14454);
	not 	XG6453 	(g16609,g14454);
	not 	XG6454 	(g16631,g14454);
	not 	XG6455 	(g17242,g14454);
	not 	XG6456 	(g17216,g14454);
	not 	XG6457 	(g16750,g14454);
	not 	XG6458 	(g17411,g14454);
	not 	XG6459 	(g16530,g14454);
	not 	XG6460 	(g16320,g14454);
	not 	XG6461 	(g16726,g14454);
	not 	XG6462 	(g17366,g14454);
	not 	XG6463 	(g16727,g14454);
	not 	XG6464 	(g17301,g14454);
	not 	XG6465 	(g16695,g14454);
	not 	XG6466 	(g16661,g14454);
	not 	XG6467 	(g16632,g14454);
	not 	XG6468 	(g17470,g14454);
	not 	XG6469 	(I18469,g13809);
	not 	XG6470 	(I17125,g13809);
	not 	XG6471 	(I17198,g13809);
	not 	XG6472 	(I18842,g13809);
	not 	XG6473 	(I17111,g13809);
	not 	XG6474 	(I18265,g13350);
	not 	XG6475 	(I18143,g13350);
	not 	XG6476 	(I18131,g13350);
	not 	XG6477 	(I17159,g13350);
	not 	XG6478 	(I18120,g13350);
	not 	XG6479 	(I17228,g13350);
	not 	XG6480 	(I18829,g13350);
	not 	XG6481 	(I18382,g13350);
	not 	XG6482 	(I18313,g13350);
	not 	XG6483 	(g17157,g13350);
	not 	XG6484 	(I17639,g13350);
	not 	XG6485 	(I18078,g13350);
	not 	XG6486 	(g17794,g13350);
	not 	XG6487 	(I18482,g13350);
	not 	XG6488 	(g17489,g12955);
	not 	XG6489 	(g17465,g12955);
	not 	XG6490 	(g17410,g12955);
	not 	XG6491 	(I17136,g14398);
	not 	XG6492 	(I18865,g14314);
	not 	XG6493 	(I17723,g13177);
	not 	XG6494 	(I18154,g13177);
	not 	XG6495 	(I18104,g13177);
	not 	XG6496 	(I18252,g13177);
	not 	XG6497 	(I18165,g13177);
	not 	XG6498 	(I17675,g13394);
	not 	XG6499 	(I17401,g13394);
	not 	XG6500 	(I17488,g13394);
	not 	XG6501 	(I17471,g13394);
	not 	XG6502 	(I18083,g13394);
	not 	XG6503 	(I17658,g13394);
	not 	XG6504 	(I17420,g13394);
	not 	XG6505 	(I17661,g13329);
	not 	XG6506 	(I18849,g14290);
	not 	XG6507 	(I17590,g14591);
	not 	XG6508 	(I17355,g14591);
	not 	XG6509 	(I17098,g14336);
	not 	XG6510 	(I17374,g13638);
	not 	XG6511 	(I17976,g13638);
	not 	XG6512 	(I18028,g13638);
	not 	XG6513 	(I18048,g13638);
	not 	XG6514 	(I18285,g13638);
	not 	XG6515 	(I17442,g13638);
	not 	XG6516 	(I18003,g13638);
	not 	XG6517 	(I18006,g13638);
	not 	XG6518 	(I18839,g13716);
	not 	XG6519 	(I18852,g13716);
	not 	XG6520 	(I18810,g13716);
	not 	XG6521 	(I18350,g13716);
	not 	XG6522 	(I17173,g13716);
	not 	XG6523 	(I17679,g13416);
	not 	XG6524 	(I17425,g13416);
	not 	XG6525 	(I17436,g13416);
	not 	XG6526 	(I18101,g13416);
	not 	XG6527 	(I17699,g13416);
	not 	XG6528 	(I17491,g13416);
	not 	XG6529 	(I17507,g13416);
	not 	XG6530 	(I17154,g13605);
	not 	XG6531 	(I17276,g13605);
	not 	XG6532 	(I18180,g13605);
	not 	XG6533 	(I17249,g13605);
	not 	XG6534 	(I18221,g13605);
	not 	XG6535 	(I18320,g13605);
	not 	XG6536 	(g17512,g12983);
	not 	XG6537 	(g17491,g12983);
	not 	XG6538 	(g17466,g12983);
	not 	XG6539 	(I17188,g13782);
	not 	XG6540 	(I18832,g13782);
	not 	XG6541 	(I18434,g13782);
	not 	XG6542 	(I17108,g13782);
	not 	XG6543 	(I18875,g13782);
	not 	XG6544 	(I18868,g14315);
	not 	XG6545 	(I17704,g13144);
	not 	XG6546 	(I18089,g13144);
	not 	XG6547 	(I18151,g13144);
	not 	XG6548 	(I18135,g13144);
	not 	XG6549 	(I18238,g13144);
	not 	XG6550 	(I17101,g14338);
	not 	XG6551 	(I17104,g12932);
	not 	XG6552 	(I18855,g13745);
	not 	XG6553 	(I18398,g13745);
	not 	XG6554 	(I18822,g13745);
	not 	XG6555 	(I17181,g13745);
	not 	XG6556 	(I18872,g13745);
	not 	XG6557 	(I17392,g13680);
	not 	XG6558 	(I18071,g13680);
	not 	XG6559 	(I18009,g13680);
	not 	XG6560 	(I17456,g13680);
	not 	XG6561 	(I18031,g13680);
	not 	XG6562 	(I18323,g13680);
	not 	XG6563 	(I18051,g13680);
	not 	XG6564 	(I18034,g13680);
	not 	XG6565 	(I17121,g14366);
	not 	XG6566 	(I18858,g13835);
	not 	XG6567 	(I17128,g13835);
	not 	XG6568 	(I18518,g13835);
	not 	XG6569 	(I17140,g13835);
	not 	XG6570 	(I17207,g13835);
	and 	XG6571 	(g15858,g14045,g3542);
	and 	XG6572 	(g16868,g14297,g5813);
	not 	XG6573 	(g17087,g14321);
	not 	XG6574 	(g17147,g14321);
	not 	XG6575 	(g17121,g14321);
	not 	XG6576 	(g17789,g14321);
	and 	XG6577 	(g16163,g14179,g14254);
	nand 	XG6578 	(I17447,I17446,g13336);
	nand 	XG6579 	(I17884,I17883,g13336);
	nand 	XG6580 	(I17475,I17474,g13336);
	nand 	XG6581 	(I17380,I17379,g13336);
	and 	XG6582 	(g15613,g13555,g3490);
	nand 	XG6583 	(g12351,I15195,I15194);
	nor 	XG6584 	(g19209,g11320,g15614,g12971);
	nand 	XG6585 	(g17736,g12563,g5659,g14522,g5563);
	nand 	XG6586 	(g12301,I15149,I15148);
	nand 	XG6587 	(g15735,g9864,g5659,g14425,g5547);
	nand 	XG6588 	(g20172,g8131,g16876);
	nand 	XG6589 	(g20163,g13938,g16663);
	nor 	XG6590 	(g12970,g10488,g10510,g10555);
	not 	XG6591 	(g10544,I13906);
	not 	XG6592 	(g16958,g14238);
	not 	XG6593 	(g17085,g14238);
	not 	XG6594 	(g16968,g14238);
	not 	XG6595 	(g17733,g14238);
	not 	XG6596 	(g13138,I15765);
	nand 	XG6597 	(g17605,g12563,g5630,g14425,g5559);
	and 	XG6598 	(g16023,g13584,g3813);
	nand 	XG6599 	(g16815,g11631,g4005,g13824,g3909);
	nand 	XG6600 	(g15674,g13110,g921);
	and 	XG6601 	(g17783,g13110,g7851);
	or 	XG6602 	(g19356,g14874,g17784);
	nand 	XG6603 	(g17755,g9864,g5630,g14522,g5619);
	not 	XG6604 	(I16724,g12108);
	not 	XG6605 	(I16698,g12077);
	nand 	XG6606 	(g19965,g16424,g3380);
	not 	XG6607 	(I16855,g10473);
	not 	XG6608 	(g13279,I15843);
	and 	XG6609 	(g16732,g14882,g5555);
	not 	XG6610 	(g15969,I17416);
	and 	XG6611 	(g21188,g15705,g7666);
	nand 	XG6612 	(g16694,g11631,g3976,g13772,g3905);
	nand 	XG6613 	(I20467,g16728,g16663);
	nand 	XG6614 	(g12423,I15243,I15242);
	not 	XG6615 	(g16688,g14045);
	not 	XG6616 	(g16654,g14136);
	not 	XG6617 	(g16812,g13555);
	not 	XG6618 	(g16124,g13555);
	not 	XG6619 	(g16158,g13555);
	not 	XG6620 	(g16186,g13555);
	nand 	XG6621 	(I14213,I14211,g9295);
	not 	XG6622 	(g13251,I15814);
	nand 	XG6623 	(g20186,g8177,g16926);
	nand 	XG6624 	(g17679,g12563,g5681,g14425,g5611);
	and 	XG6625 	(g14185,g11744,g8686);
	and 	XG6626 	(g14221,g11823,g8686);
	nand 	XG6627 	(g16854,g8595,g3976,g13824,g3965);
	nor 	XG6628 	(g19853,g1052,g15746);
	not 	XG6629 	(g13304,I15872);
	not 	XG6630 	(g16651,g14005);
	not 	XG6631 	(g16622,g14104);
	nand 	XG6632 	(g19611,g15995,g1199,g1070);
	nand 	XG6633 	(g13057,g11294,g969);
	and 	XG6634 	(g14207,g11793,g8639);
	and 	XG6635 	(g14233,g11855,g8639);
	nor 	XG6636 	(g16024,g11890,g14216);
	nand 	XG6637 	(I17476,I17474,g1105);
	or 	XG6638 	(g17511,I18452,g11976,g14365,g14396);
	not 	XG6639 	(g14536,I16651);
	and 	XG6640 	(g15785,g14107,g3558);
	nand 	XG6641 	(I20486,g16757,g16696);
	nand 	XG6642 	(I14532,I14530,g8873);
	nand 	XG6643 	(I14531,I14530,g8840);
	and 	XG6644 	(g15672,g13458,g433);
	and 	XG6645 	(g16204,g14348,g6537);
	and 	XG6646 	(g16668,g14962,g5543);
	and 	XG6647 	(g17768,g10741,g13325);
	nand 	XG6648 	(I15168,I15166,g9823);
	and 	XG6649 	(g15978,g14032,g246);
	not 	XG6650 	(I16629,g11987);
	nand 	XG6651 	(I15167,I15166,g9904);
	nor 	XG6652 	(g17175,g13545,g1216);
	nor 	XG6653 	(g16183,g13545,g9223);
	nand 	XG6654 	(g17514,g8595,g4019,g13772,g3917);
	nand 	XG6655 	(g16956,g11631,g4019,g13824,g3925);
	not 	XG6656 	(g14031,I16289);
	not 	XG6657 	(g17086,g14297);
	not 	XG6658 	(g17014,g14297);
	not 	XG6659 	(g17772,g14297);
	not 	XG6660 	(g17135,g14297);
	nand 	XG6661 	(g17814,g12563,g5673,g14522,g5579);
	nand 	XG6662 	(g17670,g8595,g4005,g13772,g3893);
	and 	XG6663 	(g14316,g11920,g2370);
	not 	XG6664 	(g14412,I16564);
	not 	XG6665 	(g13311,I15878);
	not 	XG6666 	(g14571,I16688);
	not 	XG6667 	(g14543,I16660);
	not 	XG6668 	(g14423,I16579);
	not 	XG6669 	(g13096,I15727);
	not 	XG6670 	(g14544,I16663);
	not 	XG6671 	(g14453,I16610);
	not 	XG6672 	(g13514,I15987);
	not 	XG6673 	(g13460,I15942);
	not 	XG6674 	(g13431,I15932);
	not 	XG6675 	(g13409,I15918);
	not 	XG6676 	(g13477,I15954);
	not 	XG6677 	(g13410,I15921);
	not 	XG6678 	(g13583,I16028);
	not 	XG6679 	(g14563,I16676);
	not 	XG6680 	(g16200,g13584);
	not 	XG6681 	(g16853,g13584);
	not 	XG6682 	(g16159,g13584);
	not 	XG6683 	(g16172,g13584);
	nand 	XG6684 	(g11389,I14400,I14399);
	not 	XG6685 	(g13258,I15821);
	and 	XG6686 	(g17785,g10762,g13341);
	not 	XG6687 	(I16775,g12183);
	not 	XG6688 	(g14308,I16471);
	and 	XG6689 	(g15936,g13999,g475);
	nand 	XG6690 	(g13256,g11812,g11294,g11846);
	or 	XG6691 	(g13211,g7567,g11294);
	and 	XG6692 	(I18762,g11498,g6767,g13156);
	and 	XG6693 	(I18785,g11498,g6767,g13156);
	and 	XG6694 	(I17542,g6756,g6767,g13156);
	and 	XG6695 	(I18713,g6756,g6767,g13156);
	not 	XG6696 	(g13250,I15811);
	not 	XG6697 	(g16685,g14038);
	not 	XG6698 	(g16423,g14066);
	or 	XG6699 	(g17264,g14309,g7118);
	and 	XG6700 	(g20131,g14309,g15170);
	nand 	XG6701 	(g11350,I14370,I14369);
	and 	XG6702 	(g15693,g13474,g269);
	and 	XG6703 	(g15902,g13975,g441);
	not 	XG6704 	(g21430,g15608);
	or 	XG6705 	(g19576,g14202,g17138);
	nand 	XG6706 	(I18682,I18680,g14752);
	not 	XG6707 	(g17641,g14845);
	not 	XG6708 	(g17602,g14962);
	not 	XG6709 	(g14332,I16492);
	nand 	XG6710 	(g16264,g13223,g9158,g518);
	not 	XG6711 	(g17599,g14794);
	not 	XG6712 	(g17308,g14876);
	not 	XG6713 	(g10521,I13889);
	not 	XG6714 	(I19802,g15727);
	and 	XG6715 	(g16845,g15011,g6593);
	not 	XG6716 	(I15494,g10385);
	not 	XG6717 	(g13280,I15846);
	and 	XG6718 	(g16846,g11185,g12591,g14034);
	nand 	XG6719 	(g15713,g9864,g5673,g14425,g5571);
	not 	XG6720 	(I16590,g11966);
	nor 	XG6721 	(g20854,g17243,g5381);
	nand 	XG6722 	(g15725,g9864,g5681,g14522,g5603);
	and 	XG6723 	(g16128,g14166,g14333);
	not 	XG6724 	(g19369,g15995);
	and 	XG6725 	(g15507,g13305,g10970);
	and 	XG6726 	(g16026,g14065,g854);
	not 	XG6727 	(g14424,g11136);
	not 	XG6728 	(g14753,g11317);
	nand 	XG6729 	(I18635,I18633,g14713);
	nor 	XG6730 	(g19793,g1404,g16292);
	not 	XG6731 	(g14384,I16538);
	not 	XG6732 	(g14616,I16733);
	not 	XG6733 	(g12940,g11744);
	not 	XG6734 	(g12997,g11826);
	not 	XG6735 	(g13016,g11878);
	not 	XG6736 	(g12968,g11793);
	and 	XG6737 	(g16207,g14204,g9839);
	not 	XG6738 	(g18088,g13267);
	not 	XG6739 	(I18879,g13267);
	not 	XG6740 	(g16579,g13267);
	not 	XG6741 	(I17744,g14912);
	and 	XG6742 	(g16222,g14348,g6513);
	not 	XG6743 	(g20237,g17213);
	nor 	XG6744 	(g16210,g4894,g13479);
	and 	XG6745 	(g15863,g13223,g13762);
	and 	XG6746 	(I18620,g11498,g11450,g13156);
	and 	XG6747 	(I18765,g11498,g11450,g13156);
	and 	XG6748 	(I17741,g11498,g11450,g14988);
	and 	XG6749 	(I17552,g11498,g11450,g13156);
	and 	XG6750 	(I18819,g11498,g11450,g13156);
	and 	XG6751 	(I18740,g11498,g11450,g13156);
	and 	XG6752 	(I18568,g11498,g11450,g13156);
	and 	XG6753 	(I17585,g11498,g11450,g14988);
	and 	XG6754 	(I18671,g6756,g11450,g13156);
	and 	XG6755 	(I17529,g6756,g11450,g13156);
	and 	XG6756 	(I17606,g6756,g11450,g14988);
	and 	XG6757 	(I17575,g6756,g11450,g13156);
	and 	XG6758 	(I18782,g6756,g11450,g13156);
	and 	XG6759 	(I18716,g6756,g11450,g13156);
	and 	XG6760 	(I18803,g6756,g11450,g13156);
	and 	XG6761 	(I17692,g6756,g11450,g14988);
	or 	XG6762 	(g17464,I18385,g11935,g14313,g14334);
	not 	XG6763 	(g14307,I16468);
	not 	XG6764 	(I16515,g12477);
	not 	XG6765 	(g13271,I15834);
	not 	XG6766 	(g21510,g15647);
	not 	XG6767 	(g13024,g11900);
	not 	XG6768 	(g12998,g11829);
	not 	XG6769 	(g19533,g16261);
	not 	XG6770 	(g14443,I16596);
	and 	XG6771 	(g15852,g13223,g13820);
	and 	XG6772 	(g15903,g13223,g13796);
	and 	XG6773 	(g15876,g13223,g13512);
	not 	XG6774 	(g17616,g14309);
	not 	XG6775 	(g15811,g13125);
	not 	XG6776 	(g15799,g13110);
	not 	XG6777 	(g13007,g11852);
	not 	XG6778 	(g13015,g11875);
	not 	XG6779 	(g13033,g11917);
	not 	XG6780 	(g13045,g11941);
	not 	XG6781 	(g20070,g16173);
	and 	XG6782 	(g15745,g13223,g686);
	not 	XG6783 	(g17677,g14882);
	not 	XG6784 	(g17392,g14924);
	and 	XG6785 	(g14206,g11790,g8655);
	not 	XG6786 	(I15572,g10499);
	not 	XG6787 	(g13793,I16120);
	not 	XG6788 	(g12967,g11790);
	not 	XG6789 	(g13023,g11897);
	not 	XG6790 	(g13034,g11920);
	not 	XG6791 	(g12996,g11823);
	not 	XG6792 	(g13022,g11894);
	not 	XG6793 	(g13014,g11872);
	not 	XG6794 	(g12995,g11820);
	not 	XG6795 	(g13008,g11855);
	nor 	XG6796 	(g16479,g12490,g14719);
	not 	XG6797 	(g13510,I15981);
	or 	XG6798 	(g19522,g14180,g17057);
	not 	XG6799 	(g19427,g16292);
	not 	XG6800 	(g13303,I15869);
	nand 	XG6801 	(I14499,I14497,g8737);
	and 	XG6802 	(g16807,g14978,g6585);
	not 	XG6803 	(I16544,g11931);
	not 	XG6804 	(I16626,g11986);
	and 	XG6805 	(g16929,g14348,g6505);
	not 	XG6806 	(g21556,g15669);
	not 	XG6807 	(I16679,g12039);
	not 	XG6808 	(g17720,g15045);
	not 	XG6809 	(g17745,g14978);
	not 	XG6810 	(g17136,g14348);
	not 	XG6811 	(g17122,g14348);
	not 	XG6812 	(g17815,g14348);
	not 	XG6813 	(g17154,g14348);
	or 	XG6814 	(g17569,I18492,g11995,g14394,g14416);
	not 	XG6815 	(I16455,g11845);
	nand 	XG6816 	(I17461,I17460,g13378);
	or 	XG6817 	(g17490,I18421,g11958,g14337,g14364);
	nor 	XG6818 	(g16215,g13545,g1211);
	nor 	XG6819 	(g16226,g13545,g8052);
	not 	XG6820 	(g14358,I16512);
	not 	XG6821 	(I18370,g14873);
	nand 	XG6822 	(g20645,g17243,g14344);
	nand 	XG6823 	(I17448,I17446,g956);
	nand 	XG6824 	(g20870,g9567,g17315,g14432);
	not 	XG6825 	(g17763,g15011);
	not 	XG6826 	(g17507,g15030);
	not 	XG6827 	(g13857,I16163);
	nor 	XG6828 	(g16227,g13574,g1554);
	nor 	XG6829 	(g16237,g13574,g8088);
	not 	XG6830 	(g20085,g16187);
	not 	XG6831 	(g14442,I16593);
	not 	XG6832 	(g16325,g13223);
	not 	XG6833 	(g16712,g13223);
	not 	XG6834 	(g16289,g13223);
	not 	XG6835 	(g16680,g13223);
	not 	XG6836 	(g16310,g13223);
	not 	XG6837 	(g16768,g13223);
	not 	XG6838 	(g16739,g13223);
	and 	XG6839 	(g15873,g14072,g3550);
	not 	XG6840 	(I16541,g11929);
	nor 	XG6841 	(g17180,g13574,g1559);
	nor 	XG6842 	(g16198,g13574,g9247);
	not 	XG6843 	(g13298,I15862);
	not 	XG6844 	(g13064,g11705);
	not 	XG6845 	(g16721,g14072);
	not 	XG6846 	(g16475,g14107);
	not 	XG6847 	(I16969,g13943);
	not 	XG6848 	(g14331,I16489);
	not 	XG6849 	(I16160,g11237);
	and 	XG6850 	(g16098,g14238,g5148);
	and 	XG6851 	(g15847,g14005,g3191);
	not 	XG6852 	(I17324,g14119);
	not 	XG6853 	(I17733,g14844);
	not 	XG6854 	(I17302,g14044);
	not 	XG6855 	(I17772,g14888);
	not 	XG6856 	(I17801,g14936);
	not 	XG6857 	(I17873,g15017);
	not 	XG6858 	(I17314,g14078);
	not 	XG6859 	(I17834,g14977);
	and 	XG6860 	(g15633,g13584,g3841);
	and 	XG6861 	(g15836,g14104,g3187);
	and 	XG6862 	(g16177,g14238,g5128);
	nand 	XG6863 	(g16097,g10998,g13319);
	nand 	XG6864 	(g19530,g10841,g15829);
	and 	XG6865 	(g19350,g13505,g15968);
	and 	XG6866 	(g15701,g13584,g3821);
	and 	XG6867 	(g15874,g14079,g3893);
	nand 	XG6868 	(g13476,g11869,g11336,g7503);
	nand 	XG6869 	(g13496,g11815,g11336,g1351);
	nand 	XG6870 	(g13130,g11336,g11815,g1351);
	nand 	XG6871 	(g13554,g1351,g7582,g11336);
	and 	XG6872 	(g15653,g13530,g3119);
	and 	XG6873 	(g16161,g14297,g5841);
	nand 	XG6874 	(I18538,I18536,g14642);
	and 	XG6875 	(g16666,g14794,g5200);
	and 	XG6876 	(g21333,g15740,g1300);
	nand 	XG6877 	(I17462,I17460,g1300);
	and 	XG6878 	(g15589,g13334,g411);
	and 	XG6879 	(g14256,g11872,g2079);
	and 	XG6880 	(g16203,g14297,g5821);
	and 	XG6881 	(g16733,g14889,g5893);
	and 	XG6882 	(g14257,g11878,g8612);
	and 	XG6883 	(g14220,g11820,g8612);
	and 	XG6884 	(g16125,g14238,g5152);
	nand 	XG6885 	(I18487,I18485,g14611);
	nand 	XG6886 	(g16687,g11519,g3325,g13700,g3255);
	and 	XG6887 	(g15654,g13584,g3845);
	or 	XG6888 	(g17488,I18417,g11954,g14335,g14361);
	and 	XG6889 	(g13252,g699,g11469,g11511,g11561);
	nor 	XG6890 	(g15718,g11330,g13858);
	nor 	XG6891 	(g17515,g10828,g13221);
	and 	XG6892 	(g15757,g14066,g3207);
	nor 	XG6893 	(g16220,g4939,g13499);
	and 	XG6894 	(g16178,g14297,g5845);
	and 	XG6895 	(g15857,g14038,g3199);
	nand 	XG6896 	(g19614,g16047,g1542);
	and 	XG6897 	(g16765,g15045,g6581);
	nor 	XG6898 	(g19932,g16296,g3376);
	and 	XG6899 	(g16599,g15030,g6601);
	and 	XG6900 	(g14295,g11894,g1811);
	and 	XG6901 	(g16025,g14063,g446);
	nor 	XG6902 	(g15724,g11374,g13858);
	and 	XG6903 	(g16193,g14348,g6533);
	nand 	XG6904 	(g19265,g15710,g13091,g15715,g15721);
	and 	XG6905 	(g21302,g15731,g956);
	and 	XG6906 	(g15966,g13555,g3462);
	nand 	XG6907 	(g15717,g13092,g10754);
	nor 	XG6908 	(g19778,g1061,g16268);
	or 	XG6909 	(g13543,g10565,g10543);
	nand 	XG6910 	(g21253,g17482,g6423);
	or 	XG6911 	(g19336,g14831,g17769);
	nand 	XG6912 	(I17495,I17494,g13378);
	nand 	XG6913 	(I17924,I17923,g13378);
	nand 	XG6914 	(I17405,I17404,g13378);
	and 	XG6915 	(g14296,g11897,g2638);
	nand 	XG6916 	(I18681,I18680,g2638);
	or 	XG6917 	(g20187,g13491,g16202);
	or 	XG6918 	(g19587,g13046,g15700);
	and 	XG6919 	(g15567,g13312,g392);
	nand 	XG6920 	(I17381,I17379,g1129);
	and 	XG6921 	(g15673,g13437,g182);
	nand 	XG6922 	(g13079,g11336,g1312);
	nand 	XG6923 	(I14498,I14497,g9020);
	nand 	XG6924 	(g15864,g12487,g12543,g14833);
	nand 	XG6925 	(g15833,g12337,g12378,g14714);
	not 	XG6926 	(g14645,I16755);
	and 	XG6927 	(g17809,g13125,g7873);
	nand 	XG6928 	(g15695,g13125,g1266);
	nand 	XG6929 	(g15723,g13104,g10775);
	nor 	XG6930 	(g19873,g1395,g15755);
	and 	XG6931 	(g16485,g14924,g5563);
	and 	XG6932 	(g16751,g13065,g13155);
	nand 	XG6933 	(g15572,g7219,g12969);
	nand 	XG6934 	(I18634,I18633,g2504);
	nand 	XG6935 	(g13459,g11846,g11294,g7479);
	nand 	XG6936 	(g13475,g11786,g11294,g1008);
	nand 	XG6937 	(g13528,g1008,g7549,g11294);
	nand 	XG6938 	(g13115,g11294,g11786,g1008);
	or 	XG6939 	(g17510,I18449,g11972,g14362,g14393);
	and 	XG6940 	(g15651,g13414,g429);
	and 	XG6941 	(g16184,g14183,g9285);
	or 	XG6942 	(g15935,g10665,g13029);
	nand 	XG6943 	(g17598,g8595,g4027,g13824,g3949);
	and 	XG6944 	(g16806,g14971,g6247);
	and 	XG6945 	(g16701,g14845,g5547);
	nand 	XG6946 	(g19597,g15995,g1199);
	and 	XG6947 	(g20751,g4836,g16260);
	and 	XG6948 	(g14222,g11826,g8655);
	and 	XG6949 	(g16801,g14238,g5120);
	and 	XG6950 	(g21361,g16066,g7869);
	nand 	XG6951 	(g20871,g17396,g14434);
	nand 	XG6952 	(g15726,g10003,g6365,g14529,g6263);
	or 	XG6953 	(g16810,g11032,g13461);
	and 	XG6954 	(g17365,g13036,g7650);
	and 	XG6955 	(g15706,g13484,g13296);
	and 	XG6956 	(g17752,g13174,g7841);
	and 	XG6957 	(g16191,g14262,g5475);
	and 	XG6958 	(g15937,g14387,g11950);
	and 	XG6959 	(g17770,g13189,g7863);
	and 	XG6960 	(g20108,g11048,g15508);
	and 	XG6961 	(g20093,g14584,g15372);
	or 	XG6962 	(g19605,g13063,g15707);
	nand 	XG6963 	(g17820,g12614,g6019,g14549,g5925);
	nand 	XG6964 	(g20173,g13972,g16696);
	nand 	XG6965 	(g15853,g12337,g9417,g14714);
	nand 	XG6966 	(g15907,g12487,g9417,g14833);
	and 	XG6967 	(g16122,g14291,g9491);
	nand 	XG6968 	(g17297,g14291,g2729);
	nor 	XG6969 	(g16231,g4771,g13515);
	nand 	XG6970 	(g17872,g12721,g6711,g14602,g6617);
	and 	XG6971 	(g13019,g11737,g194);
	or 	XG6972 	(g19344,g14832,g17771);
	or 	XG6973 	(g18994,g13632,g16303);
	nand 	XG6974 	(g12471,I15289,I15288);
	nand 	XG6975 	(g17792,g12721,g6697,g14602,g6601);
	nand 	XG6976 	(I18589,I18587,g14679);
	not 	XG6977 	(g16206,g13437);
	not 	XG6978 	(g16235,g13437);
	not 	XG6979 	(g16214,g13437);
	not 	XG6980 	(g17056,g13437);
	not 	XG6981 	(g16195,g13437);
	not 	XG6982 	(g16223,g13437);
	not 	XG6983 	(g16180,g13437);
	not 	XG6984 	(g16127,g13437);
	not 	XG6985 	(g16162,g13437);
	not 	XG6986 	(g16099,g13437);
	not 	XG6987 	(I18233,g14639);
	nor 	XG6988 	(g16646,g11372,g11020,g13437);
	nand 	XG6989 	(I18581,I18579,g14678);
	nand 	XG6990 	(I18580,I18579,g1945);
	or 	XG6991 	(g19501,g14168,g16986);
	nor 	XG6992 	(g16201,g4704,g13462);
	not 	XG6993 	(g16966,g14291);
	nand 	XG6994 	(g16770,g8481,g3274,g13765,g3263);
	and 	XG6995 	(g19911,g17748,g14707);
	nor 	XG6996 	(g21389,g12259,g17748,g10143);
	nand 	XG6997 	(g21190,g17420,g6077);
	not 	XG6998 	(I18148,g13526);
	and 	XG6999 	(g15849,g14136,g3538);
	and 	XG7000 	(g20875,g4681,g16281);
	nand 	XG7001 	(g20838,g17284,g5041);
	nand 	XG7002 	(g17513,g8481,g3325,g13765,g3247);
	not 	XG7003 	(g17717,g14937);
	not 	XG7004 	(g17481,g15005);
	and 	XG7005 	(g16840,g14262,g5467);
	or 	XG7006 	(g19467,g14097,g16896);
	nor 	XG7007 	(g16219,g4760,g13498);
	nand 	XG7008 	(g16625,g11519,g3274,g13700,g3203);
	not 	XG7009 	(I21162,g17292);
	and 	XG7010 	(g16633,g14921,g5196);
	nand 	XG7011 	(g17846,g12672,g6365,g14575,g6271);
	nand 	XG7012 	(g19632,g16047,g1542,g1413);
	not 	XG7013 	(g13413,g11737);
	and 	XG7014 	(g16427,g14876,g5216);
	and 	XG7015 	(g16224,g14232,g14583);
	nand 	XG7016 	(I17406,I17404,g1472);
	and 	XG7017 	(g15679,g13555,g3470);
	not 	XG7018 	(g16514,g14139);
	not 	XG7019 	(g16724,g14079);
	or 	XG7020 	(g19274,g14791,g17753);
	and 	XG7021 	(g16735,g15027,g6235);
	not 	XG7022 	(g17120,g14262);
	not 	XG7023 	(g17754,g14262);
	not 	XG7024 	(g17013,g14262);
	not 	XG7025 	(g16969,g14262);
	nor 	XG7026 	(g16232,g4950,g13516);
	nand 	XG7027 	(g17734,g9780,g5283,g14490,g5272);
	nand 	XG7028 	(g17578,g12497,g5283,g14399,g5212);
	or 	XG7029 	(g19557,g14190,g17123);
	or 	XG7030 	(g20202,g13507,g16211);
	nand 	XG7031 	(g16749,g11631,g4027,g13772,g3957);
	or 	XG7032 	(g19488,g14148,g16965);
	or 	XG7033 	(g19619,g13080,g15712);
	nand 	XG7034 	(g15709,g9780,g5327,g14399,g5224);
	nand 	XG7035 	(g16741,g11519,g3303,g13765,g3207);
	nand 	XG7036 	(g17597,g8481,g3303,g13700,g3191);
	not 	XG7037 	(g17419,g14965);
	not 	XG7038 	(g17680,g14889);
	or 	XG7039 	(g19595,g14218,g17149);
	nand 	XG7040 	(I14332,I14330,g9966);
	not 	XG7041 	(g20272,g17239);
	not 	XG7042 	(g16691,g14160);
	not 	XG7043 	(g16747,g14113);
	or 	XG7044 	(g20217,g13523,g16221);
	not 	XG7045 	(g21413,g15585);
	and 	XG7046 	(g21378,g16090,g7887);
	not 	XG7047 	(g19518,g16239);
	and 	XG7048 	(g21298,g15825,g7697);
	nand 	XG7049 	(g19506,g15825,g4087);
	or 	XG7050 	(g13242,g7601,g11336);
	nand 	XG7051 	(g13264,g11849,g11336,g11869);
	nand 	XG7052 	(I18588,I18587,g2370);
	nand 	XG7053 	(I17496,I17494,g1448);
	nand 	XG7054 	(g11419,I14429,I14428);
	and 	XG7055 	(g16212,g14321,g6167);
	not 	XG7056 	(g21460,g15628);
	and 	XG7057 	(g16700,g14838,g5208);
	not 	XG7058 	(g17644,g15002);
	not 	XG7059 	(g17714,g14930);
	nand 	XG7060 	(I14331,I14330,g225);
	or 	XG7061 	(g19475,g14126,g16930);
	nand 	XG7062 	(g17765,g12721,g6719,g14556,g6649);
	and 	XG7063 	(g15590,g13530,g3139);
	nor 	XG7064 	(g16287,g11144,g13622);
	and 	XG7065 	(g19275,g16044,g7823);
	not 	XG7066 	(I19762,g15732);
	and 	XG7067 	(g16884,g14321,g6159);
	and 	XG7068 	(g21285,g16027,g7857);
	and 	XG7069 	(g16192,g14321,g6191);
	and 	XG7070 	(g16179,g14321,g6187);
	not 	XG7071 	(g16171,g13530);
	not 	XG7072 	(g16096,g13530);
	not 	XG7073 	(g16769,g13530);
	not 	XG7074 	(g16123,g13530);
	or 	XG7075 	(g20276,g13566,g16243);
	not 	XG7076 	(g19407,g16268);
	and 	XG7077 	(g15632,g13555,g3494);
	nand 	XG7078 	(g19857,g16296,g13628);
	or 	XG7079 	(g19879,g13265,g15841);
	nand 	XG7080 	(I14212,I14211,g9252);
	and 	XG7081 	(g21296,g16072,g7879);
	nand 	XG7082 	(g15753,g10003,g6351,g14529,g6239);
	nand 	XG7083 	(g17640,g12497,g5335,g14399,g5264);
	or 	XG7084 	(g19363,g14913,g17810);
	not 	XG7085 	(g19362,g16072);
	not 	XG7086 	(g19428,g16090);
	or 	XG7087 	(g19604,g13059,g15704);
	nand 	XG7088 	(g12239,I15107,I15106);
	nand 	XG7089 	(g17708,g12497,g5313,g14490,g5216);
	nand 	XG7090 	(g17775,g12672,g6351,g14575,g6255);
	not 	XG7091 	(g19364,g15825);
	or 	XG7092 	(g20241,g13541,g16233);
	and 	XG7093 	(g19207,g15992,g7803);
	nand 	XG7094 	(I17885,I17883,g1135);
	and 	XG7095 	(g20887,g4864,g16282);
	nand 	XG7096 	(g17790,g10003,g6322,g14575,g6311);
	nand 	XG7097 	(g17686,g12672,g6322,g14529,g6251);
	not 	XG7098 	(g19071,g15591);
	or 	XG7099 	(g17268,g14387,g9220);
	not 	XG7100 	(g19355,g16027);
	not 	XG7101 	(g19738,g15992);
	not 	XG7102 	(g19408,g16066);
	not 	XG7103 	(g20765,g17748);
	not 	XG7104 	(g17575,g14921);
	not 	XG7105 	(g17638,g14838);
	and 	XG7106 	(g21347,g15750,g1339);
	not 	XG7107 	(g19374,g16047);
	nand 	XG7108 	(g20734,g17312,g14408);
	nand 	XG7109 	(I18537,I18536,g2236);
	not 	XG7110 	(g16809,g14387);
	not 	XG7111 	(g17683,g15027);
	not 	XG7112 	(g17742,g14971);
	not 	XG7113 	(g20212,g17194);
	nand 	XG7114 	(g21011,g9629,g17399,g14504);
	and 	XG7115 	(g15703,g13437,g452);
	and 	XG7116 	(g15722,g13437,g464);
	nand 	XG7117 	(g17635,g8542,g3654,g13730,g3542);
	nand 	XG7118 	(g17788,g12497,g5327,g14490,g5232);
	nand 	XG7119 	(g17757,g12614,g6005,g14549,g5909);
	and 	XG7120 	(g16520,g14965,g5909);
	nand 	XG7121 	(g16657,g11576,g3625,g13730,g3554);
	nand 	XG7122 	(g15729,g9935,g6027,g14549,g5949);
	nand 	XG7123 	(g17716,g12614,g6027,g14497,g5957);
	nand 	XG7124 	(g15743,g9935,g6005,g14497,g5893);
	nand 	XG7125 	(g16813,g8542,g3625,g13799,g3614);
	nor 	XG7126 	(g21140,g17312,g6073);
	nand 	XG7127 	(g15736,g10003,g6373,g14575,g6295);
	nand 	XG7128 	(g17744,g12672,g6373,g14529,g6303);
	nand 	XG7129 	(g17572,g8542,g3676,g13799,g3598);
	nand 	XG7130 	(g16875,g11519,g3317,g13765,g3223);
	nand 	XG7131 	(g17468,g8481,g3317,g13700,g3215);
	and 	XG7132 	(g15797,g14139,g3909);
	nand 	XG7133 	(g17647,g12614,g5976,g14497,g5905);
	or 	XG7134 	(g19525,g16811,g7696);
	and 	XG7135 	(g21163,g4878,g16321);
	nand 	XG7136 	(g16723,g11576,g3676,g13730,g3606);
	and 	XG7137 	(g20739,g4674,g16259);
	and 	XG7138 	(g15911,g13530,g3111);
	nor 	XG7139 	(g16488,g13656,g13697);
	and 	XG7140 	(g16538,g15005,g6255);
	and 	XG7141 	(g17636,g13463,g10829);
	and 	XG7142 	(g17671,g13485,g7685);
	and 	XG7143 	(g21024,g4871,g16306);
	nand 	XG7144 	(g17816,g10061,g6668,g14602,g6657);
	nand 	XG7145 	(g17723,g12721,g6668,g14556,g6597);
	nand 	XG7146 	(g15728,g9780,g5313,g14399,g5200);
	or 	XG7147 	(g19359,g14875,g17786);
	nand 	XG7148 	(g17773,g9935,g5976,g14549,g5965);
	or 	XG7149 	(g17594,I18543,g12025,g14420,g14450);
	and 	XG7150 	(g15612,g13530,g3143);
	nand 	XG7151 	(g17495,g8542,g3668,g13730,g3566);
	nor 	XG7152 	(g16242,g4961,g13529);
	and 	XG7153 	(g16762,g14930,g5901);
	and 	XG7154 	(g17145,g13249,g7469);
	nor 	XG7155 	(g16209,g4749,g13478);
	and 	XG7156 	(g16703,g15002,g5889);
	or 	XG7157 	(g17570,I18495,g11999,g14397,g14419);
	nand 	XG7158 	(g15719,g9780,g5335,g14490,g5256);
	nand 	XG7159 	(g20675,g9442,g17246,g14377);
	and 	XG7160 	(g15652,g13437,g174);
	nand 	XG7161 	(g16772,g11576,g3654,g13799,g3558);
	and 	XG7162 	(g16160,g14262,g5499);
	and 	XG7163 	(g15884,g14113,g3901);
	nand 	XG7164 	(g16925,g11576,g3668,g13799,g3574);
	not 	XG7165 	(g19751,g16044);
	and 	XG7166 	(g19791,g17189,g14253);
	and 	XG7167 	(g15860,g14160,g3889);
	nand 	XG7168 	(g15702,g7293,g13066);
	nor 	XG7169 	(g20717,g17217,g5037);
	and 	XG7170 	(g16126,g14262,g5495);
	nand 	XG7171 	(g15720,g9935,g6019,g14497,g5917);
	nand 	XG7172 	(g20733,g9509,g17290,g14406);
	and 	XG7173 	(g15694,g13437,g457);
	and 	XG7174 	(g15611,g13437,g471);
	and 	XG7175 	(g16763,g14937,g6239);
	nand 	XG7176 	(g19903,g8227,g16319,g13707);
	nand 	XG7177 	(g20979,g17309,g5385);
	nand 	XG7178 	(g19916,g16313,g3029);
	and 	XG7179 	(g15631,g13437,g168);
	nand 	XG7180 	(g19874,g8163,g16299,g13665);
	nor 	XG7181 	(g19887,g16275,g3025);
	and 	XG7182 	(g21332,g15739,g996);
	nand 	XG7183 	(g15581,g12999,g7232);
	nand 	XG7184 	(g15744,g10061,g6719,g14602,g6641);
	and 	XG7185 	(g15716,g13437,g468);
	and 	XG7186 	(g21012,g4688,g16304);
	and 	XG7187 	(g15711,g13437,g460);
	nand 	XG7188 	(g20676,g17287,g14379);
	nand 	XG7189 	(g15708,g13083,g7340);
	nand 	XG7190 	(g20644,g9372,g17220,g14342);
	nand 	XG7191 	(g19795,g16275,g13600);
	nand 	XG7192 	(g19875,g16316,g13667);
	nor 	XG7193 	(g21250,g17494,g9340,g9417);
	nor 	XG7194 	(g21277,g17467,g9340,g9417);
	nand 	XG7195 	(g15962,g9340,g9417,g14833);
	nand 	XG7196 	(g15877,g12543,g9340,g14833);
	nand 	XG7197 	(g15867,g9340,g9417,g14714);
	nand 	XG7198 	(g15844,g12378,g9340,g14714);
	and 	XG7199 	(g20559,g15831,g336);
	nand 	XG7200 	(I17925,I17923,g1478);
	and 	XG7201 	(g20682,g4646,g16238);
	nand 	XG7202 	(g15782,g10061,g6697,g14556,g6585);
	nand 	XG7203 	(g19856,g8105,g16278,g13626);
	nand 	XG7204 	(g15730,g10061,g6711,g14556,g6609);
	nor 	XG7205 	(g21206,g17396,g6419);
	and 	XG7206 	(g17133,g13222,g10683);
	nand 	XG7207 	(I18531,I18529,g14640);
	and 	XG7208 	(g16855,g13107,g4392);
	nand 	XG7209 	(g21124,g17393,g5731);
	nor 	XG7210 	(g17625,g12123,g14541);
	not 	XG7211 	(g20035,g16430);
	nand 	XG7212 	(I18486,I18485,g1677);
	nand 	XG7213 	(g20011,g16476,g3731);
	and 	XG7214 	(g18935,g15574,g4322);
	nand 	XG7215 	(I18627,I18625,g14712);
	not 	XG7216 	(g21306,g15582);
	nand 	XG7217 	(g20619,g17217,g14317);
	not 	XG7218 	(g19146,g15574);
	nand 	XG7219 	(I18626,I18625,g2079);
	nor 	XG7220 	(g19981,g16316,g3727);
	nor 	XG7221 	(g20995,g17287,g5727);
	nand 	XG7222 	(I18530,I18529,g1811);
	not 	XG7223 	(g15680,I17207);
	not 	XG7224 	(g15563,I17140);
	not 	XG7225 	(g17587,I18518);
	not 	XG7226 	(g15483,I17128);
	not 	XG7227 	(g17952,I18858);
	not 	XG7228 	(g15426,I17121);
	not 	XG7229 	(g16826,I18034);
	not 	XG7230 	(g16861,I18051);
	not 	XG7231 	(g17384,I18323);
	not 	XG7232 	(g16821,I18031);
	not 	XG7233 	(g16077,I17456);
	not 	XG7234 	(g16795,I18009);
	not 	XG7235 	(g16877,I18071);
	not 	XG7236 	(g15915,I17392);
	not 	XG7237 	(g18062,I18872);
	not 	XG7238 	(g15615,I17181);
	not 	XG7239 	(g17818,I18822);
	not 	XG7240 	(g17475,I18398);
	not 	XG7241 	(g17929,I18855);
	not 	XG7242 	(g15277,I17104);
	not 	XG7243 	(g15224,I17101);
	not 	XG7244 	(g17200,I18238);
	not 	XG7245 	(g16987,I18135);
	not 	XG7246 	(g17059,I18151);
	not 	XG7247 	(g16923,I18089);
	not 	XG7248 	(g16508,I17704);
	not 	XG7249 	(g18008,I18868);
	not 	XG7250 	(g18065,I18875);
	not 	XG7251 	(g15345,I17108);
	not 	XG7252 	(g17501,I18434);
	not 	XG7253 	(g17844,I18832);
	not 	XG7254 	(g15634,I17188);
	not 	XG7255 	(g17367,I18320);
	not 	XG7256 	(g17183,I18221);
	not 	XG7257 	(g15733,I17249);
	not 	XG7258 	(g17128,I18180);
	not 	XG7259 	(g15758,I17276);
	not 	XG7260 	(g15573,I17154);
	not 	XG7261 	(g16164,I17507);
	not 	XG7262 	(g16136,I17491);
	not 	XG7263 	(g16489,I17699);
	not 	XG7264 	(g16931,I18101);
	not 	XG7265 	(g16031,I17436);
	not 	XG7266 	(g16000,I17425);
	not 	XG7267 	(g16449,I17679);
	not 	XG7268 	(g15595,I17173);
	not 	XG7269 	(g17413,I18350);
	not 	XG7270 	(g17812,I18810);
	not 	XG7271 	(g17926,I18852);
	not 	XG7272 	(g17847,I18839);
	not 	XG7273 	(g16782,I18006);
	not 	XG7274 	(g16777,I18003);
	not 	XG7275 	(g16053,I17442);
	not 	XG7276 	(g17302,I18285);
	not 	XG7277 	(g16856,I18048);
	not 	XG7278 	(g16816,I18028);
	not 	XG7279 	(g16752,I17976);
	not 	XG7280 	(g15885,I17374);
	not 	XG7281 	(g15171,I17098);
	not 	XG7282 	(g15862,I17355);
	not 	XG7283 	(g16249,I17590);
	not 	XG7284 	(g17873,I18849);
	not 	XG7285 	(g16349,I17661);
	not 	XG7286 	(g15979,I17420);
	not 	XG7287 	(g16326,I17658);
	not 	XG7288 	(g16897,I18083);
	not 	XG7289 	(g16100,I17471);
	not 	XG7290 	(g16129,I17488);
	not 	XG7291 	(g15938,I17401);
	not 	XG7292 	(g16431,I17675);
	not 	XG7293 	(g17093,I18165);
	not 	XG7294 	(g17226,I18252);
	not 	XG7295 	(g16954,I18104);
	not 	XG7296 	(g17062,I18154);
	not 	XG7297 	(g16525,I17723);
	not 	XG7298 	(g17955,I18865);
	not 	XG7299 	(g15509,I17136);
	not 	XG7300 	(g17533,I18482);
	not 	XG7301 	(g16886,I18078);
	not 	XG7302 	(g16309,I17639);
	not 	XG7303 	(g17328,I18313);
	not 	XG7304 	(g17433,I18382);
	not 	XG7305 	(g17821,I18829);
	not 	XG7306 	(g15714,I17228);
	not 	XG7307 	(g16964,I18120);
	not 	XG7308 	(g15579,I17159);
	not 	XG7309 	(g16971,I18131);
	not 	XG7310 	(g17015,I18143);
	not 	XG7311 	(g17249,I18265);
	not 	XG7312 	(g15348,I17111);
	not 	XG7313 	(g17870,I18842);
	not 	XG7314 	(g15656,I17198);
	not 	XG7315 	(g15480,I17125);
	not 	XG7316 	(g17526,I18469);
	not 	XG7317 	(g16587,I17763);
	not 	XG7318 	(g16967,I18125);
	not 	XG7319 	(g17271,I18270);
	not 	XG7320 	(g17125,I18177);
	not 	XG7321 	(g17096,I18168);
	not 	XG7322 	(g15373,I17118);
	not 	XG7323 	(g15085,I17008);
	not 	XG7324 	(I18900,g16767);
	not 	XG7325 	(I18903,g16872);
	not 	XG7326 	(I18909,g16873);
	not 	XG7327 	(I18897,g16738);
	not 	XG7328 	(I18888,g16644);
	not 	XG7329 	(I18891,g16676);
	not 	XG7330 	(I18894,g16708);
	not 	XG7331 	(I18906,g16963);
	not 	XG7332 	(I18885,g16643);
	not 	XG7333 	(I18882,g16580);
	not 	XG7334 	(g17485,I18408);
	not 	XG7335 	(g17614,I18571);
	not 	XG7336 	(g17326,I18307);
	not 	XG7337 	(g17508,I18443);
	not 	XG7338 	(g17428,I18367);
	not 	XG7339 	(g16308,I17636);
	not 	XG7340 	(g17532,I18479);
	not 	XG7341 	(g17427,I18364);
	not 	XG7342 	(g16487,I17695);
	not 	XG7343 	(g17247,I18259);
	not 	XG7344 	(g17691,I18674);
	not 	XG7345 	(g16578,I17750);
	not 	XG7346 	(g17486,I18411);
	not 	XG7347 	(g16323,I17653);
	not 	XG7348 	(g17327,I18310);
	not 	XG7349 	(g17432,I18379);
	not 	XG7350 	(g17409,I18344);
	not 	XG7351 	(g17591,I18526);
	not 	XG7352 	(g17296,I18280);
	not 	XG7353 	(g17430,I18373);
	not 	XG7354 	(g17615,I18574);
	not 	XG7355 	(g17224,I18248);
	not 	XG7356 	(g17509,I18446);
	not 	XG7357 	(g17178,I18214);
	not 	XG7358 	(g17324,I18301);
	nor 	XG7359 	(g21652,g17663,g17619);
	not 	XG7360 	(g21653,g17663);
	not 	XG7361 	(I20929,g17663);
	not 	XG7362 	(I19012,g15060);
	not 	XG7363 	(I19235,g15078);
	nor 	XG7364 	(g21655,g17700,g17657);
	not 	XG7365 	(I20891,g17700);
	not 	XG7366 	(g21656,g17700);
	not 	XG7367 	(g21654,g17619);
	not 	XG7368 	(I20882,g17619);
	not 	XG7369 	(I19348,g15084);
	not 	XG7370 	(I19487,g15125);
	not 	XG7371 	(I19238,g15079);
	not 	XG7372 	(I18912,g15050);
	nor 	XG7373 	(g21658,g17727,g17694);
	not 	XG7374 	(g21660,g17694);
	not 	XG7375 	(I20793,g17694);
	not 	XG7376 	(g21659,g17727);
	not 	XG7377 	(I20840,g17727);
	not 	XG7378 	(I20830,g17657);
	not 	XG7379 	(g21657,g17657);
	not 	XG7380 	(I19345,g15083);
	not 	XG7381 	(I19484,g15122);
	not 	XG7382 	(g13856,I16160);
	not 	XG7383 	(I17094,g14331);
	not 	XG7384 	(g15048,I16969);
	and 	XG7385 	(g19393,g16325,g691);
	and 	XG7386 	(g19788,g17216,g9983);
	and 	XG7387 	(g19691,g17085,g9614);
	and 	XG7388 	(g19461,g16846,g11708);
	and 	XG7389 	(g19145,g16200,g8450);
	and 	XG7390 	(g16662,g14753,g4552);
	nand 	XG7391 	(g13241,g10544,g7503);
	nand 	XG7392 	(g13580,g10544,g7922,g7503,g11849);
	nand 	XG7393 	(g13573,g1351,g7582,g10544,g8002);
	nand 	XG7394 	(g19589,g10884,g10841,g15969);
	nand 	XG7395 	(g19546,g10884,g10841,g15969);
	nand 	XG7396 	(g19483,g10922,g10841,g15969);
	nand 	XG7397 	(g19513,g10922,g10841,g15969);
	nand 	XG7398 	(g16093,I17462,I17461);
	not 	XG7399 	(I17747,g13298);
	and 	XG7400 	(g18910,g16075,g16227);
	and 	XG7401 	(g18933,g13597,g16237);
	and 	XG7402 	(g19735,g17135,g9740);
	not 	XG7403 	(g14385,I16541);
	and 	XG7404 	(g16279,g14424,g4512);
	nand 	XG7405 	(g20783,g17225,g14616);
	and 	XG7406 	(g19717,g17122,g6527);
	and 	XG7407 	(g19736,g17136,g12136);
	nand 	XG7408 	(g20181,g16846,g13252);
	nand 	XG7409 	(g22709,g19611,g1193);
	nand 	XG7410 	(g21272,g17157,g11268);
	and 	XG7411 	(g19948,g16320,g17515);
	and 	XG7412 	(g17690,I18671,g11640,g11592,g11547);
	and 	XG7413 	(g17724,I18713,g11640,g11592,g11547);
	and 	XG7414 	(g17613,I18568,g11640,g11592,g11547);
	and 	XG7415 	(g17766,I18762,g11640,g11592,g6772);
	and 	XG7416 	(g17747,I18740,g11640,g11592,g6772);
	and 	XG7417 	(g17780,I18782,g11640,g11592,g6772);
	and 	XG7418 	(g21251,g17470,g13969);
	not 	XG7419 	(I17148,g14442);
	and 	XG7420 	(g19637,g16958,g5142);
	and 	XG7421 	(g19660,g16968,g12001);
	nand 	XG7422 	(g13918,g11350,g3267,g11217,g3259);
	nand 	XG7423 	(g19442,g17794,g11431);
	and 	XG7424 	(g19588,g16853,g3849);
	and 	XG7425 	(g20094,g16631,g8872);
	not 	XG7426 	(I18262,g13857);
	nand 	XG7427 	(g13240,g10521,g1046);
	and 	XG7428 	(g20188,g17772,g5849);
	nand 	XG7429 	(g16069,I17448,I17447);
	and 	XG7430 	(g23392,g21430,g7247);
	not 	XG7431 	(g23391,g20645);
	not 	XG7432 	(g17429,I18370);
	nand 	XG7433 	(g20784,g17595,g14616);
	and 	XG7434 	(g17140,g12968,g8616);
	and 	XG7435 	(g17176,g13008,g8616);
	not 	XG7436 	(I17114,g14358);
	nand 	XG7437 	(g21294,g17157,g11324);
	nand 	XG7438 	(g17699,I18682,I18681);
	not 	XG7439 	(g14277,I16455);
	and 	XG7440 	(g17192,g13022,g1677);
	not 	XG7441 	(g14564,I16679);
	and 	XG7442 	(g19564,g13976,g17175);
	and 	XG7443 	(g19578,g11130,g16183);
	or 	XG7444 	(g19441,g12931,g15507);
	nand 	XG7445 	(g15904,I17381,I17380);
	not 	XG7446 	(g14509,I16626);
	nand 	XG7447 	(g13058,g1312,g10544);
	not 	XG7448 	(g14386,I16544);
	nand 	XG7449 	(g11545,I14499,I14498);
	and 	XG7450 	(g20162,g16750,g8737);
	and 	XG7451 	(g21405,g15811,g13377);
	not 	XG7452 	(I17780,g13303);
	and 	XG7453 	(g19693,g17087,g6181);
	and 	XG7454 	(g19716,g17121,g12100);
	and 	XG7455 	(g20171,g10476,g16479);
	and 	XG7456 	(g20215,g10476,g16479);
	not 	XG7457 	(I17609,g13510);
	and 	XG7458 	(g17193,g13023,g2504);
	nand 	XG7459 	(g17662,I18635,I18634);
	nand 	XG7460 	(g13551,g10521,g7903,g7479,g11812);
	nand 	XG7461 	(g13210,g10521,g7479);
	nand 	XG7462 	(g15832,g13256,g7479,g7903);
	nand 	XG7463 	(g16181,g13459,g13057,g13495,g13475);
	nand 	XG7464 	(g13544,g1008,g7549,g10521,g7972);
	or 	XG7465 	(g19555,g13030,g15672);
	nand 	XG7466 	(g21403,g17157,g11652);
	nor 	XG7467 	(g19063,g15674,g7909);
	and 	XG7468 	(g21557,g15674,g12980);
	or 	XG7469 	(g20169,g13460,g16184);
	not 	XG7470 	(I18224,g13793);
	and 	XG7471 	(g18951,g16124,g3484);
	and 	XG7472 	(g18981,g16158,g11206);
	nand 	XG7473 	(g20107,g17794,g11404);
	not 	XG7474 	(g12952,I15572);
	nand 	XG7475 	(g21288,g17492,g14616);
	and 	XG7476 	(g20375,g16846,g671);
	nand 	XG7477 	(g20092,g17794,g11373);
	or 	XG7478 	(g18879,g14423,g17365);
	nand 	XG7479 	(g19510,g10899,g10841,g15969);
	nand 	XG7480 	(g19549,g10899,g10841,g15969);
	nand 	XG7481 	(g19455,g7781,g10841,g15969);
	nand 	XG7482 	(g19495,g7781,g10841,g15969);
	or 	XG7483 	(g19267,g17768,g17752);
	nand 	XG7484 	(g19886,g17794,g11403);
	nand 	XG7485 	(g21388,g17157,g11608);
	or 	XG7486 	(g20160,g13415,g16163);
	or 	XG7487 	(g19337,g17785,g17770);
	and 	XG7488 	(g18906,g16264,g13568);
	not 	XG7489 	(I18523,g14443);
	nand 	XG7490 	(g21377,g17157,g11560);
	nand 	XG7491 	(I20488,I20486,g16757);
	nor 	XG7492 	(g19907,g13676,g16210);
	nand 	XG7493 	(g21354,g17157,g11468);
	not 	XG7494 	(I17650,g13271);
	not 	XG7495 	(g14359,I16515);
	and 	XG7496 	(g20165,g17733,g5156);
	nand 	XG7497 	(g21301,g17157,g11371);
	not 	XG7498 	(I18861,g14307);
	nand 	XG7499 	(g20081,g17794,g11325);
	nand 	XG7500 	(g21331,g17157,g11402);
	not 	XG7501 	(g16540,I17744);
	not 	XG7502 	(g20033,g16579);
	not 	XG7503 	(g18091,I18879);
	not 	XG7504 	(I19917,g18088);
	not 	XG7505 	(I17131,g14384);
	nand 	XG7506 	(g21344,g17157,g11428);
	nor 	XG7507 	(g22983,g19853,g16268,g979);
	or 	XG7508 	(g20148,g13393,g16128);
	nor 	XG7509 	(g23626,g20854,g17309);
	nand 	XG7510 	(g19450,g17794,g11471);
	not 	XG7511 	(g14441,I16590);
	not 	XG7512 	(g20065,g16846);
	not 	XG7513 	(g20078,g16846);
	not 	XG7514 	(I17671,g13280);
	not 	XG7515 	(g12875,I15494);
	not 	XG7516 	(g19264,I19802);
	nand 	XG7517 	(I20468,I20467,g16663);
	not 	XG7518 	(g19609,g16264);
	and 	XG7519 	(g19069,g16186,g8397);
	nor 	XG7520 	(g23079,g19965,g8390);
	not 	XG7521 	(I18376,g14332);
	nand 	XG7522 	(g21359,g17157,g11509);
	and 	XG7523 	(g19571,g16812,g3498);
	nand 	XG7524 	(g20199,g13907,g16749,g13968,g16815);
	and 	XG7525 	(g17781,I18785,g6789,g11592,g6772);
	or 	XG7526 	(g20051,g13306,g15936);
	not 	XG7527 	(g13877,g11350);
	not 	XG7528 	(g21393,g17264);
	not 	XG7529 	(I17612,g13250);
	not 	XG7530 	(g15571,g13211);
	or 	XG7531 	(g20063,g13313,g15978);
	nand 	XG7532 	(g21353,g17157,g11467);
	not 	XG7533 	(I18341,g14308);
	not 	XG7534 	(g14676,I16775);
	not 	XG7535 	(I17633,g13258);
	not 	XG7536 	(g13902,g11389);
	not 	XG7537 	(I18205,g14563);
	not 	XG7538 	(I17808,g13311);
	not 	XG7539 	(I17143,g14412);
	and 	XG7540 	(g19746,g17147,g9816);
	not 	XG7541 	(I18476,g14031);
	nand 	XG7542 	(g12332,I15168,I15167);
	not 	XG7543 	(g14510,I16629);
	nand 	XG7544 	(g21360,g17157,g11510);
	nand 	XG7545 	(g20007,g17794,g11512);
	nand 	XG7546 	(g14739,g12351,g5983,g12067,g5929);
	and 	XG7547 	(g20977,g17301,g10123);
	nand 	XG7548 	(g11591,I14532,I14531);
	and 	XG7549 	(g20095,g16632,g8873);
	not 	XG7550 	(I17166,g14536);
	nand 	XG7551 	(g16119,I17476,I17475);
	not 	XG7552 	(I17783,g13304);
	and 	XG7553 	(g20135,g16695,g16258);
	nand 	XG7554 	(g13257,g10544,g1389);
	and 	XG7555 	(g23292,g16726,g19879);
	not 	XG7556 	(I17615,g13251);
	nand 	XG7557 	(g11154,I14213,I14212);
	not 	XG7558 	(g14745,g12423);
	nand 	XG7559 	(g19913,g17794,g11430);
	nand 	XG7560 	(g21385,g14636,g17679,g14696,g17736);
	nand 	XG7561 	(g21283,g17157,g11291);
	nand 	XG7562 	(I20469,I20467,g16728);
	nand 	XG7563 	(g20039,g17794,g11250);
	not 	XG7564 	(I17668,g13279);
	nand 	XG7565 	(g19474,g17794,g11609);
	not 	XG7566 	(g14790,I16855);
	nand 	XG7567 	(g16681,I17885,I17884);
	and 	XG7568 	(g20203,g17789,g6195);
	not 	XG7569 	(g14582,I16698);
	not 	XG7570 	(g14609,I16724);
	nand 	XG7571 	(g21345,g17157,g11429);
	nand 	XG7572 	(g14695,g12301,g5637,g12029,g5583);
	nand 	XG7573 	(g17712,g12301,g5666,g14425,g5599);
	nand 	XG7574 	(g17740,g12351,g6012,g14497,g5945);
	nand 	XG7575 	(g14771,g12351,g5969,g12129,g5961);
	not 	XG7576 	(g19502,g15674);
	nand 	XG7577 	(g21417,g17157,g11677);
	nand 	XG7578 	(g21330,g17157,g11401);
	nand 	XG7579 	(g20055,g17794,g11269);
	and 	XG7580 	(g20112,g16661,g13540);
	not 	XG7581 	(I18788,g13138);
	nand 	XG7582 	(g14730,g12301,g5623,g12093,g5615);
	nand 	XG7583 	(g20068,g17794,g11293);
	not 	XG7584 	(g14669,g12301);
	not 	XG7585 	(g14701,g12351);
	nand 	XG7586 	(g19962,g17794,g11470);
	nand 	XG7587 	(g19466,g17794,g11562);
	and 	XG7588 	(g19752,g15864,g2771);
	and 	XG7589 	(g17150,g12995,g8579);
	and 	XG7590 	(g17182,g13016,g8579);
	nand 	XG7591 	(g21287,g17571,g14616);
	nand 	XG7592 	(g16719,g11350,g3310,g13700,g3243);
	and 	XG7593 	(g19139,g16195,g452);
	and 	XG7594 	(g19333,g16223,g464);
	and 	XG7595 	(g19462,g16646,g14177,g14182,g7850);
	or 	XG7596 	(g20082,g13321,g16026);
	nand 	XG7597 	(g17593,I18538,I18537);
	and 	XG7598 	(g17199,g13034,g2236);
	and 	XG7599 	(g22859,g20734,g9456);
	and 	XG7600 	(g23412,g21510,g7297);
	not 	XG7601 	(g23411,g20734);
	nand 	XG7602 	(g21357,g13086,g15726,g13109,g15736);
	nand 	XG7603 	(g21416,g14706,g17744,g14781,g17775);
	or 	XG7604 	(g15800,g13242,g10821);
	and 	XG7605 	(g17191,g13242,g1384);
	or 	XG7606 	(g22304,g17693,g21347);
	nand 	XG7607 	(g20170,g13866,g16687,g13897,g16741);
	nand 	XG7608 	(g20111,g14422,g17468,g14517,g17513);
	and 	XG7609 	(g23229,g4521,g18994);
	and 	XG7610 	(g23151,g7162,g18994);
	nand 	XG7611 	(g13958,g11389,g3618,g11238,g3610);
	nand 	XG7612 	(g17761,g12423,g6358,g14529,g6291);
	and 	XG7613 	(g21394,g15799,g13335);
	not 	XG7614 	(g20192,g17268);
	nand 	XG7615 	(g14820,g12423,g6315,g12173,g6307);
	not 	XG7616 	(g23055,g20887);
	not 	XG7617 	(g22870,g20887);
	not 	XG7618 	(g22718,g20887);
	not 	XG7619 	(g23285,g20887);
	nand 	XG7620 	(g23132,g19932,g8155);
	or 	XG7621 	(g22152,g17469,g21188);
	nand 	XG7622 	(g23733,g11178,g20751);
	nand 	XG7623 	(g21363,g14598,g17640,g14664,g17708);
	not 	XG7624 	(g14631,g12239);
	nand 	XG7625 	(g13993,g11419,g3969,g11255,g3961);
	nand 	XG7626 	(g16776,g11419,g4012,g13772,g3945);
	nand 	XG7627 	(g14780,g12423,g6329,g12101,g6275);
	and 	XG7628 	(g19692,g17086,g12066);
	and 	XG7629 	(g19681,g17014,g5835);
	and 	XG7630 	(g22760,g20237,g9360);
	not 	XG7631 	(g22759,g19857);
	nand 	XG7632 	(g16745,g11389,g3661,g13730,g3594);
	nand 	XG7633 	(g21334,g17596,g14616);
	or 	XG7634 	(g20077,g13320,g16025);
	or 	XG7635 	(g20034,g13299,g15902);
	and 	XG7636 	(g18950,g16123,g11193);
	and 	XG7637 	(g18993,g16172,g11224);
	and 	XG7638 	(g18982,g16159,g3835);
	or 	XG7639 	(g20905,g17264,g7216);
	and 	XG7640 	(g20193,g17264,g15578);
	nand 	XG7641 	(g13043,g969,g10521);
	nand 	XG7642 	(g21187,g17364,g14616);
	nand 	XG7643 	(g17779,g12471,g6704,g14556,g6637);
	and 	XG7644 	(g18974,g16127,g174);
	and 	XG7645 	(g19914,g15853,g2815);
	and 	XG7646 	(g17151,g12996,g8659);
	and 	XG7647 	(g17091,g12940,g8659);
	nand 	XG7648 	(g21289,g17493,g14616);
	nand 	XG7649 	(g13967,g11419,g3983,g11225,g3929);
	nand 	XG7650 	(I20487,I20486,g16696);
	not 	XG7651 	(g19061,I19762);
	and 	XG7652 	(g19740,g15907,g2783);
	and 	XG7653 	(g17139,g12967,g8635);
	and 	XG7654 	(g17152,g12997,g8635);
	nand 	XG7655 	(g21186,g17363,g14616);
	or 	XG7656 	(g19575,g13042,g15693);
	or 	XG7657 	(g22226,g17655,g21333);
	nand 	XG7658 	(g19358,g1399,g15723);
	nand 	XG7659 	(g21339,g13050,g15713,g13084,g15725);
	nand 	XG7660 	(g20151,g14519,g17514,g14570,g17598);
	and 	XG7661 	(g19266,g16214,g246);
	nor 	XG7662 	(g20000,g16264,g13661);
	and 	XG7663 	(g16234,I17575,g11640,g6782,g6772);
	and 	XG7664 	(g17817,I18819,g11640,g6782,g11547);
	and 	XG7665 	(g16539,I17741,g6789,g6782,g11547);
	and 	XG7666 	(g16194,I17529,g11640,g6782,g11547);
	and 	XG7667 	(g16205,I17542,g11640,g6782,g11547);
	and 	XG7668 	(g16213,I17552,g11640,g6782,g6772);
	nand 	XG7669 	(g21307,g13040,g15709,g13067,g15719);
	and 	XG7670 	(g18893,g16030,g16215);
	and 	XG7671 	(g18909,g13570,g16226);
	and 	XG7672 	(g19601,g11149,g16198);
	and 	XG7673 	(g19585,g14004,g17180);
	nand 	XG7674 	(g21433,g14750,g17765,g14830,g17792);
	nand 	XG7675 	(g11292,I14332,I14331);
	nand 	XG7676 	(I20460,g14187,g17515);
	not 	XG7677 	(g13933,g11419);
	nand 	XG7678 	(g16155,I17496,I17495);
	nand 	XG7679 	(g17624,I18589,I18588);
	not 	XG7680 	(g15580,g13242);
	not 	XG7681 	(g22406,g19506);
	nor 	XG7682 	(g19997,g13739,g16231);
	nor 	XG7683 	(g19880,g13634,g16201);
	nand 	XG7684 	(g23666,g11139,g20875);
	and 	XG7685 	(g19354,g16235,g471);
	and 	XG7686 	(g22340,g13522,g19605);
	and 	XG7687 	(g19516,g16097,g7824);
	and 	XG7688 	(g19521,g16739,g513);
	and 	XG7689 	(g19767,g14203,g16810);
	nand 	XG7690 	(g13927,g11389,g3632,g11207,g3578);
	or 	XG7691 	(g15789,g13211,g10819);
	and 	XG7692 	(g17179,g13211,g1041);
	nand 	XG7693 	(g23978,g12323,g21389,g572);
	and 	XG7694 	(g22534,g21389,g8766);
	nand 	XG7695 	(g23659,g20854,g9434);
	and 	XG7696 	(g20109,g17616,g17954);
	nand 	XG7697 	(g13896,g11350,g3281,g11194,g3227);
	and 	XG7698 	(g18943,g16099,g269);
	or 	XG7699 	(g19535,g13020,g15651);
	and 	XG7700 	(g17793,I18803,g6789,g11592,g6772);
	and 	XG7701 	(g16244,I17585,g6789,g11592,g11547);
	and 	XG7702 	(g16283,I17606,g6789,g11592,g11547);
	and 	XG7703 	(g17767,I18765,g6789,g11592,g6772);
	and 	XG7704 	(g16486,I17692,g6789,g11592,g6772);
	and 	XG7705 	(g17725,I18716,g6789,g11592,g11547);
	and 	XG7706 	(g17653,I18620,g6789,g11592,g11547);
	and 	XG7707 	(g19680,g17013,g12028);
	nand 	XG7708 	(g14829,g12471,g6675,g12137,g6621);
	and 	XG7709 	(g19536,g16768,g518);
	nand 	XG7710 	(g15959,I17406,I17405);
	not 	XG7711 	(I20499,g16224);
	nand 	XG7712 	(g19335,g1056,g15717);
	or 	XG7713 	(g19449,g12939,g15567);
	and 	XG7714 	(g19500,g16712,g504);
	not 	XG7715 	(g21451,I21162);
	and 	XG7716 	(g20218,g17815,g6541);
	and 	XG7717 	(g19206,g16206,g460);
	and 	XG7718 	(g22762,g20645,g9305);
	nand 	XG7719 	(g16893,g703,g13252,g10685);
	not 	XG7720 	(g22869,g20875);
	not 	XG7721 	(g23402,g20875);
	not 	XG7722 	(g23931,g20875);
	not 	XG7723 	(g23645,g20875);
	not 	XG7724 	(g17058,I18148);
	not 	XG7725 	(g23182,g21389);
	nor 	XG7726 	(g23051,g19427,g7960);
	or 	XG7727 	(g20196,g13497,g16207);
	and 	XG7728 	(g19756,g17154,g9899);
	nand 	XG7729 	(g17618,I18581,I18580);
	and 	XG7730 	(g17181,g13014,g1945);
	nand 	XG7731 	(g16713,I17925,I17924);
	nand 	XG7732 	(g14871,g12471,g6661,g12211,g6653);
	and 	XG7733 	(g19487,g16680,g499);
	not 	XG7734 	(g20540,g16646);
	not 	XG7735 	(g17197,I18233);
	not 	XG7736 	(g14786,g12471);
	not 	XG7737 	(g20388,g17297);
	not 	XG7738 	(g20531,g15907);
	not 	XG7739 	(g20782,g15853);
	and 	XG7740 	(g22871,g20871,g9523);
	and 	XG7741 	(g19384,g16310,g667);
	or 	XG7742 	(g23574,g20108,g20093);
	and 	XG7743 	(g22680,g7781,g19530);
	not 	XG7744 	(I20035,g15706);
	nor 	XG7745 	(g19953,g13712,g16220);
	and 	XG7746 	(g19372,g16289,g686);
	and 	XG7747 	(g23424,g21556,g7345);
	not 	XG7748 	(g23423,g20871);
	not 	XG7749 	(g23971,g20751);
	not 	XG7750 	(g23714,g20751);
	not 	XG7751 	(g22858,g20751);
	not 	XG7752 	(g23425,g20751);
	not 	XG7753 	(g22449,g19597);
	nor 	XG7754 	(g23711,g21253,g9892);
	nor 	XG7755 	(g22993,g19873,g16292,g1322);
	and 	XG7756 	(g21605,g15695,g13005);
	not 	XG7757 	(g19524,g15695);
	not 	XG7758 	(g20572,g15833);
	not 	XG7759 	(g20550,g15864);
	nand 	XG7760 	(g17568,I18487,I18486);
	and 	XG7761 	(g16957,g10418,g13064);
	or 	XG7762 	(g19486,g12979,g15589);
	not 	XG7763 	(g16521,g13543);
	or 	XG7764 	(g22217,g17617,g21302);
	nor 	XG7765 	(g23108,g19932,g16424);
	not 	XG7766 	(g22492,g19614);
	nand 	XG7767 	(g16196,g13476,g13079,g13513,g13496);
	not 	XG7768 	(I22024,g19350);
	not 	XG7769 	(g16640,I17834);
	not 	XG7770 	(g15816,I17314);
	not 	XG7771 	(g16675,I17873);
	not 	XG7772 	(g16615,I17801);
	not 	XG7773 	(g16594,I17772);
	not 	XG7774 	(g15806,I17302);
	not 	XG7775 	(g16533,I17733);
	not 	XG7776 	(g15824,I17324);
	nand 	XG7777 	(g20248,g14123,g14146,g17056);
	nor 	XG7778 	(g21062,g17297,g9547);
	and 	XG7779 	(g19684,g17297,g2735);
	nand 	XG7780 	(g23286,g20887,g6875);
	nand 	XG7781 	(g15843,g13264,g7503,g7922);
	and 	XG7782 	(g18992,g16171,g8341);
	nor 	XG7783 	(g23560,g20838,g9607);
	nor 	XG7784 	(g23678,g21190,g9809);
	nand 	XG7785 	(g23309,g21024,g6905);
	nand 	XG7786 	(g17656,I18627,I18626);
	and 	XG7787 	(g22191,g19875,g8119);
	and 	XG7788 	(g19784,g15877,g2775);
	nand 	XG7789 	(g23909,g20739,g7028);
	and 	XG7790 	(g22846,g20676,g9386);
	and 	XG7791 	(g21348,g17625,g10121);
	and 	XG7792 	(g21303,g17625,g10120);
	and 	XG7793 	(g23381,g21413,g7239);
	not 	XG7794 	(g23380,g20619);
	and 	XG7795 	(g22172,g19857,g8064);
	nand 	XG7796 	(g17592,I18531,I18530);
	and 	XG7797 	(g19062,g16180,g446);
	nand 	XG7798 	(g22753,g19632,g1536);
	nor 	XG7799 	(g23024,g19407,g7936);
	nor 	XG7800 	(g19140,g15695,g7939);
	and 	XG7801 	(g19768,g15833,g2803);
	nand 	XG7802 	(g23756,g21206,g9621);
	not 	XG7803 	(g22311,g18935);
	and 	XG7804 	(g23900,g19408,g1129);
	nor 	XG7805 	(g23208,g16324,g20035);
	and 	XG7806 	(g18987,g16162,g182);
	and 	XG7807 	(g19661,g16969,g5489);
	nor 	XG7808 	(g21284,g9690,g16646);
	and 	XG7809 	(g19749,g16646,g732);
	or 	XG7810 	(g19572,g14193,g17133);
	or 	XG7811 	(g19904,g14654,g17636);
	or 	XG7812 	(g19593,g14210,g17145);
	or 	XG7813 	(g19949,g14681,g17671);
	nand 	XG7814 	(g23972,g20751,g7097);
	and 	XG7815 	(g19855,g15962,g2787);
	and 	XG7816 	(g20174,g17754,g5503);
	nand 	XG7817 	(g17675,g12239,g5320,g14399,g5252);
	nor 	XG7818 	(g19999,g13742,g16232);
	and 	XG7819 	(g19715,g17120,g9679);
	and 	XG7820 	(g19594,g17268,g11913);
	and 	XG7821 	(g22161,g19071,g13202);
	nor 	XG7822 	(g23729,g21206,g17482);
	nor 	XG7823 	(g19906,g13672,g16209);
	nor 	XG7824 	(g19951,g13709,g16219);
	nor 	XG7825 	(g20027,g13779,g16242);
	nand 	XG7826 	(g23890,g20682,g7004);
	and 	XG7827 	(g19655,g16966,g2729);
	and 	XG7828 	(g19545,g16769,g3147);
	nand 	XG7829 	(g21365,g13100,g15730,g13119,g15744);
	nor 	XG7830 	(g23052,g19916,g8334);
	nand 	XG7831 	(g23932,g20875,g7051);
	and 	XG7832 	(g15650,g13413,g8362);
	nor 	XG7833 	(g23602,g20979,g9672);
	nand 	XG7834 	(g23590,g11111,g20682);
	not 	XG7835 	(g23889,g20682);
	not 	XG7836 	(g23563,g20682);
	not 	XG7837 	(I23099,g20682);
	not 	XG7838 	(g22845,g20682);
	not 	XG7839 	(g23382,g20682);
	and 	XG7840 	(g22309,g19751,g1478);
	or 	XG7841 	(g22707,g17156,g20559);
	not 	XG7842 	(g20269,g15844);
	not 	XG7843 	(g20328,g15867);
	not 	XG7844 	(g20595,g15877);
	not 	XG7845 	(g20643,g15962);
	not 	XG7846 	(I22769,g21277);
	not 	XG7847 	(I22725,g21250);
	and 	XG7848 	(g22843,g20272,g9429);
	not 	XG7849 	(g22842,g19875);
	and 	XG7850 	(g23103,g20765,g10143);
	and 	XG7851 	(g22717,g20212,g9291);
	not 	XG7852 	(g22716,g19795);
	nand 	XG7853 	(g23726,g21140,g9559);
	and 	XG7854 	(g18934,g16096,g3133);
	nand 	XG7855 	(g23623,g20717,g9364);
	and 	XG7856 	(g23401,g21460,g7262);
	not 	XG7857 	(g23400,g20676);
	nand 	XG7858 	(g14663,g12239,g5290,g12002,g5236);
	nand 	XG7859 	(g23699,g11160,g21012);
	not 	XG7860 	(g23681,g21012);
	not 	XG7861 	(g23413,g21012);
	not 	XG7862 	(g23948,g21012);
	not 	XG7863 	(g22896,g21012);
	or 	XG7864 	(g22225,g17654,g21332);
	and 	XG7865 	(g23917,g19428,g1472);
	nor 	XG7866 	(g23063,g19887,g16313);
	nor 	XG7867 	(g22654,g19506,g7733);
	and 	XG7868 	(g23854,g19506,g4093);
	nand 	XG7869 	(g23139,g10756,g21163);
	nand 	XG7870 	(g14686,g12239,g5276,g12059,g5268);
	nand 	XG7871 	(g23067,g10721,g20887);
	and 	XG7872 	(g23811,g19364,g4087);
	and 	XG7873 	(g23801,g19362,g1448);
	nand 	XG7874 	(g21351,g13069,g15720,g13098,g15729);
	nor 	XG7875 	(g23586,g20717,g17284);
	nand 	XG7876 	(g20134,g14452,g17495,g14542,g17572);
	nand 	XG7877 	(g20185,g13882,g16723,g13928,g16772);
	nand 	XG7878 	(g22306,g19071,g13202,g4616,g4584);
	or 	XG7879 	(g23405,g16245,g19791);
	or 	XG7880 	(g22669,g19525,g7763);
	and 	XG7881 	(g23779,g19355,g1105);
	nand 	XG7882 	(g23342,g21163,g6928);
	nand 	XG7883 	(g21402,g14674,g17716,g14740,g17757);
	nand 	XG7884 	(g23112,g10733,g21024);
	not 	XG7885 	(g22897,g21024);
	not 	XG7886 	(g23082,g21024);
	not 	XG7887 	(g22761,g21024);
	not 	XG7888 	(g23308,g21024);
	and 	XG7889 	(g22308,g19738,g1135);
	and 	XG7890 	(g19556,g16809,g11932);
	nand 	XG7891 	(g23630,g11123,g20739);
	not 	XG7892 	(g22857,g20739);
	not 	XG7893 	(g23908,g20739);
	not 	XG7894 	(g23605,g20739);
	not 	XG7895 	(g23393,g20739);
	not 	XG7896 	(g22919,g21163);
	not 	XG7897 	(g23341,g21163);
	not 	XG7898 	(g23127,g21163);
	not 	XG7899 	(g22844,g21163);
	nor 	XG7900 	(g23695,g21140,g17420);
	nand 	XG7901 	(g23949,g21012,g7074);
	and 	XG7902 	(g21066,g17625,g10043);
	and 	XG7903 	(g19674,g15867,g2819);
	nor 	XG7904 	(g23642,g21124,g9733);
	and 	XG7905 	(g19656,g15844,g2807);
	nor 	XG7906 	(g23124,g20011,g8443);
	and 	XG7907 	(g22720,g20619,g9253);
	and 	XG7908 	(g18890,g17625,g10158);
	and 	XG7909 	(g18949,g17625,g10183);
	nand 	XG7910 	(g23105,g19887,g8097);
	and 	XG7911 	(g21382,g17625,g10086);
	and 	XG7912 	(g22160,g19795,g8005);
	and 	XG7913 	(g21276,g17625,g10157);
	and 	XG7914 	(g21067,g17625,g10085);
	nand 	XG7915 	(g23692,g20995,g9501);
	nand 	XG7916 	(g23167,g19981,g8219);
	nor 	XG7917 	(g23662,g20995,g17393);
	nor 	XG7918 	(g23135,g19981,g16476);
	and 	XG7919 	(g18709,g17302,g59);
	and 	XG7920 	(g18374,g15171,g1878);
	and 	XG7921 	(g18282,g16136,g1379);
	and 	XG7922 	(g18343,g17955,g12847);
	and 	XG7923 	(g18420,g15373,g1996);
	and 	XG7924 	(g18671,g15758,g4628);
	and 	XG7925 	(g18656,g17128,g15120);
	nor 	XG7926 	(g19890,g8058,g16987);
	and 	XG7927 	(g18602,g16987,g3115);
	and 	XG7928 	(g18305,g16489,g1521);
	and 	XG7929 	(g18774,g15615,g5698);
	and 	XG7930 	(g18588,g16349,g2970);
	and 	XG7931 	(g18727,g16077,g4931);
	and 	XG7932 	(g18756,g15595,g5348);
	and 	XG7933 	(g18749,g17847,g5148);
	not 	XG7934 	(g18660,I19484);
	and 	XG7935 	(g18494,g15426,g2527);
	and 	XG7936 	(g18397,g15373,g2004);
	and 	XG7937 	(g18134,g17249,g534);
	and 	XG7938 	(g18161,g17433,g691);
	and 	XG7939 	(g18641,g17096,g3841);
	and 	XG7940 	(g18233,g16326,g1094);
	and 	XG7941 	(g18598,g16349,g3003);
	and 	XG7942 	(g18505,g15509,g2583);
	and 	XG7943 	(g18663,g17367,g4311);
	and 	XG7944 	(g18409,g15373,g2084);
	and 	XG7945 	(g18354,g17955,g1792);
	and 	XG7946 	(g18676,g15758,g4358);
	and 	XG7947 	(g18686,g15885,g4659);
	and 	XG7948 	(g18601,g16987,g3106);
	and 	XG7949 	(g18315,g16931,g1548);
	and 	XG7950 	(g18745,g17847,g5128);
	and 	XG7951 	(g18392,g15171,g1988);
	and 	XG7952 	(g18520,g15509,g2661);
	and 	XG7953 	(g18171,g17433,g728);
	and 	XG7954 	(g18534,g15277,g2735);
	and 	XG7955 	(g18637,g17096,g3821);
	and 	XG7956 	(g18604,g16987,g3125);
	and 	XG7957 	(g18567,g16349,g2894);
	and 	XG7958 	(g18201,g15938,g15061);
	and 	XG7959 	(g18616,g17200,g6875);
	and 	XG7960 	(g18743,g17847,g5115);
	and 	XG7961 	(g18341,g17873,g1648);
	and 	XG7962 	(g18276,g16136,g1351);
	and 	XG7963 	(g18603,g16987,g3119);
	and 	XG7964 	(g18458,g15224,g2357);
	and 	XG7965 	(g18581,g16349,g2912);
	and 	XG7966 	(g18783,g18065,g5841);
	and 	XG7967 	(g18483,g15426,g2453);
	and 	XG7968 	(g18439,g18008,g2250);
	and 	XG7969 	(g18712,g15915,g4843);
	and 	XG7970 	(g18269,g16031,g15069);
	and 	XG7971 	(g18789,g15634,g6035);
	not 	XG7972 	(g18527,I19345);
	and 	XG7973 	(g18106,g17015,g411);
	and 	XG7974 	(g18215,g15979,g943);
	and 	XG7975 	(g18307,g16931,g1559);
	and 	XG7976 	(g18633,g17226,g6905);
	and 	XG7977 	(g18698,g16777,g15131);
	and 	XG7978 	(g18410,g15373,g2079);
	and 	XG7979 	(g18779,g18065,g5821);
	and 	XG7980 	(g18612,g17200,g3329);
	nor 	XG7981 	(g19919,g11205,g16987);
	and 	XG7982 	(g18605,g16987,g3129);
	and 	XG7983 	(g18569,g16349,g94);
	and 	XG7984 	(g18659,g17183,g4366);
	and 	XG7985 	(g18406,g15373,g2060);
	and 	XG7986 	(g18274,g16031,g1311);
	and 	XG7987 	(g18230,g16326,g1111);
	and 	XG7988 	(g18582,g16349,g2922);
	and 	XG7989 	(g18540,g15277,g2775);
	and 	XG7990 	(g18757,g15595,g5352);
	nor 	XG7991 	(g20841,g12027,g17847);
	and 	XG7992 	(g18752,g17926,g15146);
	and 	XG7993 	(g18583,g16349,g2936);
	and 	XG7994 	(g18333,g17873,g1691);
	and 	XG7995 	(g18816,g15483,g6527);
	and 	XG7996 	(g18338,g17873,g1710);
	and 	XG7997 	(g18472,g15224,g2413);
	and 	XG7998 	(g18235,g16326,g1141);
	and 	XG7999 	(g18495,g15426,g2533);
	and 	XG8000 	(g18524,g15509,g2681);
	and 	XG8001 	(g18335,g17873,g1687);
	and 	XG8002 	(g18417,g15373,g2116);
	and 	XG8003 	(g18644,g17125,g15098);
	nor 	XG8004 	(g20014,g11244,g17096);
	and 	XG8005 	(g18344,g17955,g1740);
	and 	XG8006 	(g18482,g15426,g2472);
	and 	XG8007 	(g18138,g17249,g546);
	and 	XG8008 	(g18775,g15615,g7028);
	and 	XG8009 	(g18157,g17433,g15057);
	and 	XG8010 	(g18164,g17433,g699);
	and 	XG8011 	(g18454,g15224,g2303);
	and 	XG8012 	(g18593,g16349,g2999);
	and 	XG8013 	(g18362,g17955,g1834);
	and 	XG8014 	(g18212,g15979,g947);
	and 	XG8015 	(g18202,g15938,g907);
	and 	XG8016 	(g18455,g15224,g2327);
	and 	XG8017 	(g18245,g16431,g1193);
	nor 	XG8018 	(g19402,g13133,g15979);
	and 	XG8019 	(g18419,g15373,g2051);
	and 	XG8020 	(g18145,g17533,g582);
	and 	XG8021 	(g18462,g15224,g2361);
	and 	XG8022 	(g18425,g18008,g2161);
	and 	XG8023 	(g18280,g16136,g1367);
	and 	XG8024 	(g18340,g17873,g1720);
	and 	XG8025 	(g18543,g15277,g2779);
	and 	XG8026 	(g18386,g15171,g1964);
	and 	XG8027 	(g18763,g17929,g5481);
	and 	XG8028 	(g18631,g17226,g3694);
	and 	XG8029 	(g18748,g17847,g5142);
	and 	XG8030 	(g18728,g16821,g4939);
	and 	XG8031 	(g18767,g17929,g15150);
	nor 	XG8032 	(g21143,g9517,g15348);
	and 	XG8033 	(g18795,g15348,g6163);
	and 	XG8034 	(g18375,g15171,g1902);
	and 	XG8035 	(g18185,g17328,g790);
	and 	XG8036 	(g18737,g16826,g4975);
	nor 	XG8037 	(g21127,g12099,g18065);
	and 	XG8038 	(g18786,g15345,g15156);
	and 	XG8039 	(g18643,g17096,g3849);
	and 	XG8040 	(g18311,g16931,g1554);
	and 	XG8041 	(g18693,g16053,g4717);
	and 	XG8042 	(g18708,g16782,g4818);
	and 	XG8043 	(g18304,g16489,g1542);
	and 	XG8044 	(g18808,g15656,g6390);
	and 	XG8045 	(g18391,g15171,g1982);
	and 	XG8046 	(g18571,g16349,g2856);
	and 	XG8047 	(g18329,g17873,g1612);
	and 	XG8048 	(g18390,g15171,g1978);
	and 	XG8049 	(g18563,g16349,g2890);
	and 	XG8050 	(g18739,g16826,g5008);
	and 	XG8051 	(g18675,g15758,g4349);
	and 	XG8052 	(g18370,g15171,g1874);
	and 	XG8053 	(g18487,g15426,g2441);
	and 	XG8054 	(g18358,g17955,g1811);
	and 	XG8055 	(g18741,g17384,g15143);
	and 	XG8056 	(g18369,g15171,g12848);
	not 	XG8057 	(g20773,I20830);
	and 	XG8058 	(g24141,g21656,g17657);
	and 	XG8059 	(g18773,g15615,g5694);
	and 	XG8060 	(g18303,g16489,g1536);
	nor 	XG8061 	(g19422,g13141,g16031);
	and 	XG8062 	(g18691,g16053,g4727);
	and 	XG8063 	(g18817,g15483,g6533);
	and 	XG8064 	(g18278,g16136,g1345);
	and 	XG8065 	(g18584,g16349,g2950);
	and 	XG8066 	(g18302,g16489,g1514);
	and 	XG8067 	(g18131,g16971,g482);
	and 	XG8068 	(g18236,g16326,g15065);
	and 	XG8069 	(g18500,g15426,g2421);
	and 	XG8070 	(g18433,g18008,g2197);
	and 	XG8071 	(g18785,g18065,g5849);
	and 	XG8072 	(g18347,g17955,g1756);
	and 	XG8073 	(g18211,g15979,g15062);
	and 	XG8074 	(g18427,g18008,g2181);
	and 	XG8075 	(g18617,g17062,g3462);
	and 	XG8076 	(g18228,g16129,g1061);
	and 	XG8077 	(g18300,g16489,g1306);
	nor 	XG8078 	(g19338,g1306,g16031);
	and 	XG8079 	(g18824,g15680,g6732);
	and 	XG8080 	(g18411,g15373,g2093);
	and 	XG8081 	(g18327,g17873,g1636);
	and 	XG8082 	(g18165,g17433,g650);
	and 	XG8083 	(g18592,g16349,g2994);
	nor 	XG8084 	(g20720,g9299,g17847);
	and 	XG8085 	(g18744,g17847,g5124);
	and 	XG8086 	(g18268,g16000,g1280);
	and 	XG8087 	(g18489,g15426,g2509);
	and 	XG8088 	(g18361,g17955,g1821);
	and 	XG8089 	(g18558,g15277,g2803);
	and 	XG8090 	(g18266,g16000,g1274);
	and 	XG8091 	(g18121,g17015,g424);
	and 	XG8092 	(g18721,g16077,g15138);
	and 	XG8093 	(g18553,g15277,g2827);
	and 	XG8094 	(g18253,g16897,g1211);
	and 	XG8095 	(g18559,g15277,g12856);
	and 	XG8096 	(g18506,g15509,g2571);
	and 	XG8097 	(g18424,g18008,g2165);
	and 	XG8098 	(g18238,g16326,g1152);
	and 	XG8099 	(g18404,g15373,g2066);
	and 	XG8100 	(g18275,g16136,g15070);
	and 	XG8101 	(g18434,g18008,g2217);
	and 	XG8102 	(g18146,g17533,g595);
	and 	XG8103 	(g18324,g17873,g1644);
	and 	XG8104 	(g18415,g15373,g2108);
	and 	XG8105 	(g18668,g17367,g4322);
	and 	XG8106 	(g18516,g15509,g2638);
	and 	XG8107 	(g18535,g15277,g2741);
	nor 	XG8108 	(g20982,g12065,g17929);
	and 	XG8109 	(g18764,g17929,g5485);
	and 	XG8110 	(g18365,g17955,g1848);
	and 	XG8111 	(g18522,g15509,g2671);
	and 	XG8112 	(g18403,g15373,g2028);
	and 	XG8113 	(g18332,g17873,g1677);
	and 	XG8114 	(g18760,g17929,g5462);
	and 	XG8115 	(g18325,g17873,g1624);
	and 	XG8116 	(g18378,g15171,g1932);
	and 	XG8117 	(g18259,g16000,g15068);
	and 	XG8118 	(g18258,g16897,g1221);
	and 	XG8119 	(g18810,g15483,g6505);
	and 	XG8120 	(g18342,g17873,g1592);
	and 	XG8121 	(g18104,g17015,g392);
	and 	XG8122 	(g18360,g17955,g1830);
	and 	XG8123 	(g18441,g18008,g2246);
	and 	XG8124 	(g18436,g18008,g2227);
	and 	XG8125 	(g18234,g16326,g1129);
	and 	XG8126 	(g18112,g17015,g182);
	and 	XG8127 	(g18163,g17433,g79);
	and 	XG8128 	(g18160,g17433,g645);
	and 	XG8129 	(g18277,g16136,g1312);
	and 	XG8130 	(g18367,g17955,g1783);
	and 	XG8131 	(g18541,g15277,g2767);
	and 	XG8132 	(g18576,g16349,g2868);
	and 	XG8133 	(g18471,g15224,g2407);
	and 	XG8134 	(g18547,g15277,g121);
	and 	XG8135 	(g18449,g15224,g12852);
	and 	XG8136 	(g18428,g18008,g2169);
	and 	XG8137 	(g18717,g15915,g4849);
	and 	XG8138 	(g18484,g15426,g2491);
	not 	XG8139 	(g20781,I20840);
	and 	XG8140 	(g24144,g21660,g17727);
	and 	XG8141 	(g18435,g18008,g2173);
	and 	XG8142 	(g18478,g15426,g2445);
	and 	XG8143 	(g18822,g15680,g6723);
	nor 	XG8144 	(g20857,g9380,g17929);
	and 	XG8145 	(g18761,g17929,g5471);
	and 	XG8146 	(g18536,g15277,g2748);
	and 	XG8147 	(g18126,g16971,g15054);
	and 	XG8148 	(g18765,g17929,g5489);
	and 	XG8149 	(g18267,g16000,g1266);
	and 	XG8150 	(g18459,g15224,g2331);
	and 	XG8151 	(g18376,g15171,g1913);
	not 	XG8152 	(g20705,I20793);
	and 	XG8153 	(g18285,g16164,g1395);
	and 	XG8154 	(g18753,g15595,g15148);
	and 	XG8155 	(g18806,g15656,g6381);
	and 	XG8156 	(g18799,g15348,g6181);
	and 	XG8157 	(g18653,g16249,g4176);
	and 	XG8158 	(g18317,g17873,g12846);
	and 	XG8159 	(g18408,g15373,g2070);
	and 	XG8160 	(g18646,g17271,g4031);
	and 	XG8161 	(g18568,g16349,g37);
	and 	XG8162 	(g18431,g18008,g2185);
	and 	XG8163 	(g18298,g16489,g15073);
	and 	XG8164 	(g18490,g15426,g2504);
	and 	XG8165 	(g18176,g17328,g732);
	nor 	XG8166 	(g21209,g9575,g15483);
	and 	XG8167 	(g18812,g15483,g6509);
	and 	XG8168 	(g18718,g15915,g4854);
	and 	XG8169 	(g18349,g17955,g1768);
	and 	XG8170 	(g18218,g16100,g1008);
	and 	XG8171 	(g18359,g17955,g1825);
	and 	XG8172 	(g18371,g15171,g1870);
	and 	XG8173 	(g18107,g17015,g429);
	and 	XG8174 	(g18372,g15171,g1886);
	and 	XG8175 	(g18150,g17533,g604);
	and 	XG8176 	(g18412,g15373,g2098);
	and 	XG8177 	(g18210,g15938,g936);
	and 	XG8178 	(g18530,g15277,g2715);
	and 	XG8179 	(g18513,g15509,g2575);
	and 	XG8180 	(g18479,g15426,g2449);
	and 	XG8181 	(g18623,g17062,g3484);
	and 	XG8182 	(g18262,g16000,g1259);
	and 	XG8183 	(g18184,g17328,g785);
	and 	XG8184 	(g18826,g15680,g7097);
	and 	XG8185 	(g18538,g15277,g2759);
	and 	XG8186 	(g18270,g16031,g1291);
	and 	XG8187 	(g18544,g15277,g2791);
	and 	XG8188 	(g18456,g15224,g2338);
	and 	XG8189 	(g18246,g16431,g1199);
	and 	XG8190 	(g18713,g15915,g4836);
	and 	XG8191 	(g18678,g15758,g66);
	and 	XG8192 	(g18523,g15509,g2675);
	and 	XG8193 	(g18273,g16031,g1287);
	and 	XG8194 	(g18542,g15277,g2787);
	and 	XG8195 	(g18477,g15426,g2429);
	and 	XG8196 	(g18466,g15224,g2389);
	and 	XG8197 	(g18742,g17847,g5120);
	and 	XG8198 	(g18400,g15373,g2012);
	and 	XG8199 	(g18680,g15885,g15128);
	and 	XG8200 	(g18232,g16326,g1124);
	not 	XG8201 	(g18102,I18912);
	and 	XG8202 	(g18768,g17929,g5503);
	and 	XG8203 	(g18734,g16826,g4966);
	and 	XG8204 	(g18265,g16000,g1270);
	and 	XG8205 	(g18389,g15171,g1974);
	and 	XG8206 	(g18443,g18008,g2265);
	and 	XG8207 	(g18159,g17433,g671);
	and 	XG8208 	(g18260,g16000,g1252);
	and 	XG8209 	(g18162,g17433,g686);
	and 	XG8210 	(g18590,g16349,g2917);
	and 	XG8211 	(g18797,g15348,g6173);
	and 	XG8212 	(g18183,g17328,g781);
	and 	XG8213 	(g18706,g16782,g4785);
	and 	XG8214 	(g18531,g15277,g2719);
	and 	XG8215 	(g18720,g16795,g15137);
	and 	XG8216 	(g18504,g15509,g2579);
	and 	XG8217 	(g18447,g18008,g2208);
	and 	XG8218 	(g18414,g15373,g2102);
	and 	XG8219 	(g18480,g15426,g2437);
	and 	XG8220 	(g18488,g15426,g2495);
	and 	XG8221 	(g18366,g17955,g1854);
	and 	XG8222 	(g18578,g16349,g2873);
	and 	XG8223 	(g18205,g15938,g904);
	and 	XG8224 	(g18174,g17328,g739);
	and 	XG8225 	(g18762,g17929,g5475);
	and 	XG8226 	(g18147,g17533,g599);
	and 	XG8227 	(g18193,g17821,g837);
	and 	XG8228 	(g18263,g16000,g1249);
	and 	XG8229 	(g18192,g17821,g817);
	and 	XG8230 	(g18208,g15938,g930);
	and 	XG8231 	(g18158,g17433,g667);
	and 	XG8232 	(g18554,g15277,g2831);
	and 	XG8233 	(g18321,g17873,g1620);
	and 	XG8234 	(g18142,g17533,g577);
	and 	XG8235 	(g18401,g15373,g2036);
	and 	XG8236 	(g18206,g15938,g918);
	and 	XG8237 	(g18642,g17096,g15097);
	and 	XG8238 	(g18724,g16077,g4907);
	and 	XG8239 	(g18674,g15758,g4340);
	and 	XG8240 	(g18595,g16349,g2927);
	and 	XG8241 	(g18689,g16752,g15129);
	and 	XG8242 	(g18736,g16826,g4991);
	and 	XG8243 	(g18758,g15595,g7004);
	and 	XG8244 	(g18533,g15277,g2729);
	and 	XG8245 	(g18153,g17533,g626);
	and 	XG8246 	(g18529,g15277,g2712);
	and 	XG8247 	(g18444,g18008,g2269);
	and 	XG8248 	(g18615,g17200,g3347);
	and 	XG8249 	(g18609,g16987,g3147);
	and 	XG8250 	(g18701,g16856,g4771);
	and 	XG8251 	(g18445,g18008,g2273);
	and 	XG8252 	(g18792,g15634,g7051);
	and 	XG8253 	(g18387,g15171,g1955);
	and 	XG8254 	(g18256,g16897,g1242);
	and 	XG8255 	(g18751,g17847,g5156);
	and 	XG8256 	(g18501,g15509,g12854);
	and 	XG8257 	(g18295,g16449,g1489);
	and 	XG8258 	(g18515,g15509,g2643);
	and 	XG8259 	(g18492,g15426,g2523);
	and 	XG8260 	(g18364,g17955,g1844);
	and 	XG8261 	(g18152,g17533,g613);
	and 	XG8262 	(g18546,g15277,g2795);
	and 	XG8263 	(g18399,g15373,g2024);
	and 	XG8264 	(g18658,g17183,g15121);
	and 	XG8265 	(g18465,g15224,g2384);
	and 	XG8266 	(g18216,g15979,g967);
	and 	XG8267 	(g18463,g15224,g2375);
	and 	XG8268 	(g18328,g17873,g1657);
	and 	XG8269 	(g18499,g15426,g2476);
	and 	XG8270 	(g18682,g15885,g4646);
	and 	XG8271 	(g18254,g16897,g1236);
	and 	XG8272 	(g18182,g17328,g776);
	and 	XG8273 	(g18220,g16100,g1002);
	and 	XG8274 	(g18127,g16971,g499);
	and 	XG8275 	(g18719,g16795,g4894);
	and 	XG8276 	(g18572,g16349,g2864);
	nor 	XG8277 	(g19968,g11223,g17062);
	and 	XG8278 	(g18622,g17062,g3480);
	and 	XG8279 	(g18385,g15171,g1959);
	and 	XG8280 	(g18297,g16449,g1478);
	and 	XG8281 	(g18384,g15171,g1945);
	and 	XG8282 	(g18136,g17249,g550);
	and 	XG8283 	(g18448,g18008,g2153);
	and 	XG8284 	(g18497,g15426,g2541);
	and 	XG8285 	(g18725,g16077,g4912);
	and 	XG8286 	(g18549,g15277,g2799);
	and 	XG8287 	(g18379,g15171,g1906);
	and 	XG8288 	(g18248,g16897,g15067);
	and 	XG8289 	(g18574,g16349,g2882);
	and 	XG8290 	(g18813,g15483,g6513);
	and 	XG8291 	(g18306,g16931,g15074);
	and 	XG8292 	(g18151,g17533,g617);
	and 	XG8293 	(g18575,g16349,g2878);
	and 	XG8294 	(g18688,g16752,g4704);
	and 	XG8295 	(g18532,g15277,g2724);
	nor 	XG8296 	(g19984,g8171,g17096);
	and 	XG8297 	(g18636,g17096,g3817);
	and 	XG8298 	(g18286,g16164,g1404);
	and 	XG8299 	(g18320,g17873,g1616);
	and 	XG8300 	(g18591,g16349,g2965);
	and 	XG8301 	(g18791,g15634,g6044);
	and 	XG8302 	(g18141,g17533,g568);
	and 	XG8303 	(g18502,g15509,g2567);
	and 	XG8304 	(g18491,g15426,g2518);
	and 	XG8305 	(g18723,g16077,g4922);
	and 	XG8306 	(g18293,g16449,g1484);
	and 	XG8307 	(g18197,g17821,g854);
	and 	XG8308 	(g18667,g17367,g4601);
	and 	XG8309 	(g18299,g16489,g1526);
	nor 	XG8310 	(g21256,g12179,g15483);
	and 	XG8311 	(g18815,g15483,g6523);
	and 	XG8312 	(g18818,g15483,g15165);
	and 	XG8313 	(g18526,g15509,g2555);
	and 	XG8314 	(g18191,g17821,g827);
	and 	XG8315 	(g18155,g17533,g15056);
	and 	XG8316 	(g18577,g16349,g2988);
	and 	XG8317 	(g18377,g15171,g1894);
	and 	XG8318 	(g18521,g15509,g2667);
	and 	XG8319 	(g18684,g15885,g4681);
	and 	XG8320 	(g18240,g16431,g15066);
	and 	XG8321 	(g18608,g16987,g15087);
	and 	XG8322 	(g18606,g16987,g3133);
	and 	XG8323 	(g18811,g15483,g6500);
	and 	XG8324 	(g18638,g17096,g3827);
	nor 	XG8325 	(g19935,g8113,g17062);
	and 	XG8326 	(g18619,g17062,g3466);
	and 	XG8327 	(g18733,g16877,g15141);
	and 	XG8328 	(g18825,g15680,g6736);
	and 	XG8329 	(g18519,g15509,g2648);
	and 	XG8330 	(g18460,g15224,g2351);
	not 	XG8331 	(g18422,I19238);
	nor 	XG8332 	(g20998,g9450,g18065);
	and 	XG8333 	(g18778,g18065,g5817);
	and 	XG8334 	(g18692,g16053,g4732);
	and 	XG8335 	(g18679,g15758,g4633);
	and 	XG8336 	(g18654,g16249,g4146);
	and 	XG8337 	(g18405,g15373,g2040);
	and 	XG8338 	(g18196,g17821,g703);
	and 	XG8339 	(g18771,g15615,g5685);
	and 	XG8340 	(g18630,g17226,g3689);
	and 	XG8341 	(g18187,g17328,g794);
	and 	XG8342 	(g18669,g17367,g4608);
	and 	XG8343 	(g18430,g18008,g2204);
	and 	XG8344 	(g18645,g17271,g15100);
	and 	XG8345 	(g18166,g17433,g655);
	and 	XG8346 	(g18115,g17015,g460);
	and 	XG8347 	(g18759,g17929,g5467);
	not 	XG8348 	(g18661,I19487);
	and 	XG8349 	(g18363,g17955,g1840);
	and 	XG8350 	(g18699,g16816,g4760);
	and 	XG8351 	(g18330,g17873,g1668);
	and 	XG8352 	(g18819,g15483,g6541);
	and 	XG8353 	(g18398,g15373,g2020);
	and 	XG8354 	(g18467,g15224,g2380);
	and 	XG8355 	(g18685,g15885,g4688);
	and 	XG8356 	(g18780,g18065,g5827);
	and 	XG8357 	(g18125,g16886,g15053);
	and 	XG8358 	(g18452,g15224,g2311);
	and 	XG8359 	(g18509,g15509,g2587);
	and 	XG8360 	(g18128,g16971,g504);
	and 	XG8361 	(g18382,g15171,g1936);
	and 	XG8362 	(g18284,g16164,g15071);
	not 	XG8363 	(g18528,I19348);
	and 	XG8364 	(g18700,g16816,g15132);
	and 	XG8365 	(g18566,g16349,g2860);
	and 	XG8366 	(g18662,g17367,g15126);
	and 	XG8367 	(g18251,g16897,g996);
	and 	XG8368 	(g18690,g16053,g15130);
	and 	XG8369 	(g18113,g17015,g405);
	and 	XG8370 	(g18772,g15615,g5689);
	and 	XG8371 	(g18139,g17249,g542);
	and 	XG8372 	(g18292,g16449,g1472);
	and 	XG8373 	(g18508,g15509,g2606);
	and 	XG8374 	(g18137,g17249,g538);
	and 	XG8375 	(g18129,g16971,g518);
	and 	XG8376 	(g18620,g17062,g3470);
	and 	XG8377 	(g18334,g17873,g1696);
	not 	XG8378 	(g20915,I20882);
	and 	XG8379 	(g24139,g21653,g17619);
	and 	XG8380 	(g18510,g15509,g2625);
	and 	XG8381 	(g18237,g16326,g1146);
	and 	XG8382 	(g18279,g16136,g1361);
	and 	XG8383 	(g18555,g15277,g2834);
	and 	XG8384 	(g18730,g16861,g4950);
	and 	XG8385 	(g18170,g17433,g661);
	and 	XG8386 	(g18468,g15224,g2393);
	and 	XG8387 	(g18429,g18008,g2193);
	and 	XG8388 	(g18517,g15509,g2652);
	and 	XG8389 	(g18350,g17955,g1779);
	and 	XG8390 	(g18322,g17873,g1608);
	and 	XG8391 	(g18241,g16431,g1183);
	and 	XG8392 	(g18512,g15509,g2619);
	and 	XG8393 	(g18143,g17533,g586);
	and 	XG8394 	(g18626,g17062,g3498);
	and 	XG8395 	(g18446,g18008,g2279);
	and 	XG8396 	(g18351,g17955,g1760);
	and 	XG8397 	(g18635,g17096,g3808);
	and 	XG8398 	(g18110,g17015,g441);
	and 	XG8399 	(g18790,g15634,g6040);
	and 	XG8400 	(g18103,g17015,g401);
	and 	XG8401 	(g18613,g17200,g3338);
	and 	XG8402 	(g18625,g17062,g15092);
	and 	XG8403 	(g18556,g15277,g2823);
	and 	XG8404 	(g18116,g17015,g168);
	and 	XG8405 	(g18589,g16349,g2902);
	and 	XG8406 	(g18199,g17821,g832);
	and 	XG8407 	(g18189,g17821,g812);
	and 	XG8408 	(g18395,g15373,g12849);
	and 	XG8409 	(g18252,g16897,g990);
	and 	XG8410 	(g18119,g17015,g475);
	and 	XG8411 	(g18657,g17128,g4308);
	and 	XG8412 	(g18156,g17533,g572);
	and 	XG8413 	(g18514,g15509,g2629);
	and 	XG8414 	(g18373,g15171,g1890);
	and 	XG8415 	(g18696,g16053,g4741);
	and 	XG8416 	(g18353,g17955,g1772);
	and 	XG8417 	(g18475,g15426,g12853);
	not 	XG8418 	(g20922,I20891);
	and 	XG8419 	(g18611,g17200,g15090);
	and 	XG8420 	(g18801,g15348,g15160);
	and 	XG8421 	(g18135,g17249,g136);
	and 	XG8422 	(g18496,g15426,g2537);
	and 	XG8423 	(g18507,g15509,g2595);
	and 	XG8424 	(g18225,g16100,g1041);
	and 	XG8425 	(g18314,g16931,g1585);
	and 	XG8426 	(g18402,g15373,g2047);
	and 	XG8427 	(g18551,g15277,g2811);
	and 	XG8428 	(g18453,g15224,g2315);
	and 	XG8429 	(g18407,g15373,g2016);
	and 	XG8430 	(g18777,g18065,g5808);
	and 	XG8431 	(g18432,g18008,g2223);
	and 	XG8432 	(g18687,g15885,g4664);
	and 	XG8433 	(g18461,g15224,g2307);
	and 	XG8434 	(g18747,g17847,g5138);
	and 	XG8435 	(g18383,g15171,g1950);
	and 	XG8436 	(g18264,g16000,g1263);
	and 	XG8437 	(g18213,g15979,g952);
	and 	XG8438 	(g18704,g16782,g4793);
	and 	XG8439 	(g18539,g15277,g2763);
	and 	XG8440 	(g18561,g15277,g2841);
	and 	XG8441 	(g18132,g16971,g513);
	and 	XG8442 	(g18336,g17873,g1700);
	not 	XG8443 	(g18421,I19235);
	and 	XG8444 	(g18470,g15224,g2403);
	and 	XG8445 	(g18493,g15426,g2514);
	and 	XG8446 	(g18639,g17096,g3831);
	and 	XG8447 	(g18738,g16826,g15142);
	and 	XG8448 	(g18357,g17955,g1816);
	and 	XG8449 	(g18814,g15483,g6519);
	and 	XG8450 	(g18261,g16000,g1256);
	and 	XG8451 	(g18118,g17015,g471);
	and 	XG8452 	(g18537,g15277,g6856);
	and 	XG8453 	(g18120,g17015,g457);
	and 	XG8454 	(g18481,g15426,g2461);
	and 	XG8455 	(g18290,g16449,g1467);
	and 	XG8456 	(g18648,g17271,g4045);
	and 	XG8457 	(g18221,g16100,g1018);
	and 	XG8458 	(g18242,g16431,g962);
	nor 	XG8459 	(g19268,g962,g15979);
	and 	XG8460 	(g18579,g16349,g2984);
	and 	XG8461 	(g18705,g16782,g4801);
	and 	XG8462 	(g18310,g16931,g1333);
	and 	XG8463 	(g18464,g15224,g2370);
	and 	XG8464 	(g18289,g16449,g1448);
	and 	XG8465 	(g18511,g15509,g2599);
	and 	XG8466 	(g18796,g15348,g6167);
	and 	XG8467 	(g18597,g16349,g2975);
	and 	XG8468 	(g18308,g16931,g6832);
	and 	XG8469 	(g18423,g18008,g12851);
	and 	XG8470 	(g18766,g17929,g5495);
	and 	XG8471 	(g18457,g15224,g2319);
	and 	XG8472 	(g18316,g16931,g1564);
	and 	XG8473 	(g18437,g18008,g2241);
	and 	XG8474 	(g18313,g16931,g1430);
	and 	XG8475 	(g18223,g16100,g1030);
	and 	XG8476 	(g18570,g16349,g2848);
	and 	XG8477 	(g18249,g16897,g1216);
	and 	XG8478 	(g18781,g18065,g5831);
	and 	XG8479 	(g18665,g17367,g4584);
	and 	XG8480 	(g18124,g16886,g102);
	and 	XG8481 	(g18607,g16987,g3139);
	and 	XG8482 	(g18130,g16971,g528);
	and 	XG8483 	(g18707,g16782,g15134);
	and 	XG8484 	(g18672,g15758,g15127);
	and 	XG8485 	(g18649,g17271,g4049);
	and 	XG8486 	(g18250,g16897,g6821);
	and 	XG8487 	(g18326,g17873,g1664);
	and 	XG8488 	(g18621,g17062,g3476);
	not 	XG8489 	(g18200,I19012);
	and 	XG8490 	(g18820,g15563,g15166);
	and 	XG8491 	(g18677,g15758,g4639);
	and 	XG8492 	(g18651,g16249,g15102);
	and 	XG8493 	(g18178,g17328,g758);
	and 	XG8494 	(g18108,g17015,g433);
	and 	XG8495 	(g18272,g16031,g1283);
	and 	XG8496 	(g18416,g15373,g2112);
	and 	XG8497 	(g18545,g15277,g2783);
	and 	XG8498 	(g18281,g16136,g1373);
	and 	XG8499 	(g18729,g16821,g15139);
	and 	XG8500 	(g18585,g16349,g2960);
	and 	XG8501 	(g18769,g18062,g15151);
	and 	XG8502 	(g18355,g17955,g1748);
	and 	XG8503 	(g18203,g15938,g911);
	and 	XG8504 	(g18552,g15277,g2815);
	and 	XG8505 	(g18440,g18008,g2255);
	and 	XG8506 	(g18793,g15348,g6159);
	and 	XG8507 	(g18473,g15224,g2342);
	and 	XG8508 	(g18231,g16326,g1105);
	and 	XG8509 	(g18255,g16897,g1087);
	and 	XG8510 	(g18331,g17873,g1682);
	and 	XG8511 	(g18111,g17015,g174);
	and 	XG8512 	(g18629,g17226,g3680);
	and 	XG8513 	(g18803,g15480,g15161);
	nor 	XG8514 	(g21193,g12135,g15348);
	and 	XG8515 	(g18650,g17271,g6928);
	and 	XG8516 	(g18548,g15277,g2807);
	and 	XG8517 	(g18219,g16100,g969);
	and 	XG8518 	(g18754,g15595,g5339);
	and 	XG8519 	(g18204,g15938,g914);
	and 	XG8520 	(g18190,g17821,g822);
	and 	XG8521 	(g18226,g16129,g15064);
	and 	XG8522 	(g18722,g16077,g4917);
	and 	XG8523 	(g18800,g15348,g6187);
	and 	XG8524 	(g18640,g17096,g3835);
	and 	XG8525 	(g18476,g15426,g2433);
	and 	XG8526 	(g18368,g17955,g1728);
	and 	XG8527 	(g18681,g15885,g4653);
	and 	XG8528 	(g18485,g15426,g2465);
	and 	XG8529 	(g18418,g15373,g2122);
	and 	XG8530 	(g18227,g16129,g1052);
	and 	XG8531 	(g18173,g17328,g736);
	and 	XG8532 	(g18396,g15373,g2008);
	and 	XG8533 	(g18697,g16777,g4749);
	and 	XG8534 	(g18123,g16886,g479);
	and 	XG8535 	(g18807,g15656,g6386);
	and 	XG8536 	(g18784,g18065,g15155);
	and 	XG8537 	(g18318,g17873,g1604);
	and 	XG8538 	(g18627,g17093,g15093);
	and 	XG8539 	(g18586,g16349,g2886);
	and 	XG8540 	(g18109,g17015,g437);
	and 	XG8541 	(g18168,g17433,g681);
	and 	XG8542 	(g18105,g17015,g417);
	and 	XG8543 	(g18565,g16349,g2852);
	and 	XG8544 	(g18550,g15277,g2819);
	and 	XG8545 	(g18442,g18008,g2259);
	and 	XG8546 	(g18726,g16077,g4927);
	and 	XG8547 	(g18732,g16877,g4961);
	and 	XG8548 	(g18614,g17200,g3343);
	and 	XG8549 	(g18573,g16349,g2898);
	and 	XG8550 	(g18610,g17059,g15088);
	and 	XG8551 	(g18740,g17384,g4572);
	and 	XG8552 	(g18735,g16826,g4983);
	and 	XG8553 	(g18469,g15224,g2399);
	and 	XG8554 	(g18244,g16431,g1171);
	and 	XG8555 	(g18782,g18065,g5835);
	and 	XG8556 	(g18337,g17873,g1706);
	and 	XG8557 	(g18294,g16449,g15072);
	and 	XG8558 	(g18474,g15224,g2287);
	and 	XG8559 	(g18243,g16431,g1189);
	and 	XG8560 	(g18702,g16856,g15133);
	and 	XG8561 	(g18426,g18008,g2177);
	and 	XG8562 	(g18301,g16489,g1532);
	and 	XG8563 	(g18710,g17302,g15135);
	and 	XG8564 	(g18823,g15680,g6727);
	and 	XG8565 	(g18587,g16349,g2980);
	and 	XG8566 	(g18628,g17226,g15095);
	and 	XG8567 	(g18271,g16031,g1296);
	and 	XG8568 	(g18186,g17328,g753);
	and 	XG8569 	(g18288,g16449,g1454);
	and 	XG8570 	(g18770,g15615,g15153);
	and 	XG8571 	(g18525,g15509,g2610);
	and 	XG8572 	(g18673,g15758,g4643);
	and 	XG8573 	(g18287,g16449,g1442);
	and 	XG8574 	(g18695,g16053,g4737);
	and 	XG8575 	(g18175,g17328,g744);
	and 	XG8576 	(g18393,g15171,g1917);
	and 	XG8577 	(g18346,g17955,g1752);
	and 	XG8578 	(g18312,g16931,g1579);
	and 	XG8579 	(g18794,g15348,g6154);
	and 	XG8580 	(g18291,g16449,g1437);
	and 	XG8581 	(g18296,g16449,g1495);
	and 	XG8582 	(g18323,g17873,g1632);
	and 	XG8583 	(g18144,g17533,g590);
	and 	XG8584 	(g18694,g16053,g4722);
	and 	XG8585 	(g18715,g15915,g4871);
	and 	XG8586 	(g18179,g17328,g763);
	and 	XG8587 	(g18596,g16349,g2941);
	and 	XG8588 	(g18352,g17955,g1798);
	and 	XG8589 	(g18207,g15938,g925);
	and 	XG8590 	(g18486,g15426,g2485);
	and 	XG8591 	(g18746,g17847,g5134);
	and 	XG8592 	(g18172,g17328,g15058);
	and 	XG8593 	(g18133,g17249,g15055);
	and 	XG8594 	(g18755,g15595,g5343);
	and 	XG8595 	(g18809,g15656,g7074);
	and 	XG8596 	(g18239,g16326,g1135);
	and 	XG8597 	(g18802,g15348,g6195);
	and 	XG8598 	(g18167,g17433,g718);
	and 	XG8599 	(g18247,g16431,g1178);
	and 	XG8600 	(g18750,g17847,g15145);
	and 	XG8601 	(g18224,g16100,g1036);
	and 	XG8602 	(g18714,g15915,g4864);
	and 	XG8603 	(g18214,g15979,g939);
	and 	XG8604 	(g18560,g15277,g2837);
	and 	XG8605 	(g18594,g16349,g12858);
	and 	XG8606 	(g18600,g16987,g3111);
	and 	XG8607 	(g18154,g17533,g622);
	and 	XG8608 	(g18664,g17367,g4332);
	and 	XG8609 	(g18194,g17821,g843);
	and 	XG8610 	(g18169,g17433,g676);
	and 	XG8611 	(g18394,g15171,g1862);
	and 	XG8612 	(g18683,g15885,g4674);
	and 	XG8613 	(g18380,g15171,g1926);
	and 	XG8614 	(g18716,g15915,g4878);
	and 	XG8615 	(g18229,g16326,g1099);
	and 	XG8616 	(g18198,g17821,g15059);
	and 	XG8617 	(g18599,g16349,g2955);
	and 	XG8618 	(g18209,g15938,g921);
	and 	XG8619 	(g18257,g16897,g1205);
	and 	XG8620 	(g18149,g17533,g608);
	and 	XG8621 	(g18148,g17533,g562);
	and 	XG8622 	(g18634,g17096,g3813);
	and 	XG8623 	(g18787,g15634,g15158);
	and 	XG8624 	(g18731,g16861,g15140);
	and 	XG8625 	(g18413,g15373,g2089);
	and 	XG8626 	(g18804,g15656,g15163);
	and 	XG8627 	(g18180,g17328,g767);
	and 	XG8628 	(g18222,g16100,g1024);
	and 	XG8629 	(g18564,g16349,g2844);
	and 	XG8630 	(g18309,g16931,g1339);
	and 	XG8631 	(g18283,g16136,g1384);
	and 	XG8632 	(g18451,g15224,g2295);
	and 	XG8633 	(g18821,g15680,g15168);
	and 	XG8634 	(g18666,g17367,g4593);
	and 	XG8635 	(g18703,g16782,g4776);
	and 	XG8636 	(g18503,g15509,g2563);
	and 	XG8637 	(g18618,g17062,g3457);
	and 	XG8638 	(g18805,g15656,g6377);
	and 	XG8639 	(g18798,g15348,g6177);
	and 	XG8640 	(g18181,g17328,g772);
	and 	XG8641 	(g18122,g17015,g15052);
	and 	XG8642 	(g18518,g15509,g2657);
	not 	XG8643 	(g21061,I20929);
	and 	XG8644 	(g18670,g15758,g4621);
	and 	XG8645 	(g18388,g15171,g1968);
	and 	XG8646 	(g18345,g17955,g1736);
	and 	XG8647 	(g18632,g17226,g3698);
	and 	XG8648 	(g18438,g18008,g2236);
	and 	XG8649 	(g18339,g17873,g1714);
	and 	XG8650 	(g18319,g17873,g1600);
	and 	XG8651 	(g18624,g17062,g3490);
	and 	XG8652 	(g18177,g17328,g749);
	and 	XG8653 	(g18711,g15915,g15136);
	and 	XG8654 	(g18652,g16249,g4172);
	and 	XG8655 	(g18217,g16100,g15063);
	and 	XG8656 	(g18195,g17821,g847);
	and 	XG8657 	(g18788,g15634,g6031);
	and 	XG8658 	(g18188,g17328,g807);
	and 	XG8659 	(g18356,g17955,g1802);
	and 	XG8660 	(g18348,g17955,g1744);
	and 	XG8661 	(g18580,g16349,g2907);
	and 	XG8662 	(g18776,g18065,g5813);
	and 	XG8663 	(g18117,g17015,g464);
	and 	XG8664 	(g18114,g17015,g452);
	and 	XG8665 	(g18140,g17533,g559);
	and 	XG8666 	(g18498,g15426,g2547);
	and 	XG8667 	(g18647,g17271,g4040);
	and 	XG8668 	(g18450,g15224,g2299);
	and 	XG8669 	(g18381,g15171,g1882);
	and 	XG8670 	(g18557,g15277,g2771);
	not 	XG8671 	(g19638,g17324);
	not 	XG8672 	(g19417,g17178);
	not 	XG8673 	(g19376,g17509);
	not 	XG8674 	(g19757,g17224);
	not 	XG8675 	(g19773,g17615);
	not 	XG8676 	(g21222,g17430);
	not 	XG8677 	(g19620,g17296);
	not 	XG8678 	(g19345,g17591);
	not 	XG8679 	(g19626,g17409);
	not 	XG8680 	(g19662,g17432);
	not 	XG8681 	(g19379,g17327);
	not 	XG8682 	(g21370,g16323);
	not 	XG8683 	(g18984,g17486);
	not 	XG8684 	(g20204,g16578);
	not 	XG8685 	(g20097,g17691);
	not 	XG8686 	(g21156,g17247);
	not 	XG8687 	(g20277,g16487);
	not 	XG8688 	(g18954,g17427);
	not 	XG8689 	(g19389,g17532);
	not 	XG8690 	(g20242,g16308);
	not 	XG8691 	(g21225,g17428);
	not 	XG8692 	(g21160,g17508);
	not 	XG8693 	(g19330,g17326);
	not 	XG8694 	(g19606,g17614);
	not 	XG8695 	(g21308,g17485);
	not 	XG8696 	(g18093,I18885);
	not 	XG8697 	(I19384,g15085);
	not 	XG8698 	(g18876,g15373);
	not 	XG8699 	(g20503,g15373);
	not 	XG8700 	(g21408,g15373);
	not 	XG8701 	(g21274,g15373);
	not 	XG8702 	(g21422,g15373);
	not 	XG8703 	(g20609,g15373);
	not 	XG8704 	(g20664,g15373);
	not 	XG8705 	(g21179,g15373);
	not 	XG8706 	(g20914,g15373);
	not 	XG8707 	(g20665,g15373);
	not 	XG8708 	(g21054,g15373);
	not 	XG8709 	(g20704,g15373);
	not 	XG8710 	(g20383,g15373);
	not 	XG8711 	(g20444,g15373);
	not 	XG8712 	(g20545,g15373);
	not 	XG8713 	(g18887,g15373);
	not 	XG8714 	(g21052,g15373);
	not 	XG8715 	(g20634,g15373);
	not 	XG8716 	(g20564,g15373);
	not 	XG8717 	(g20663,g15373);
	not 	XG8718 	(g21454,g15373);
	not 	XG8719 	(g20913,g15373);
	not 	XG8720 	(g21053,g15373);
	not 	XG8721 	(g20703,g15373);
	not 	XG8722 	(g20587,g15373);
	not 	XG8723 	(g20502,g15373);
	not 	XG8724 	(g19800,g17096);
	not 	XG8725 	(g19677,g17096);
	not 	XG8726 	(g19861,g17096);
	not 	XG8727 	(g20238,g17096);
	not 	XG8728 	(g19771,g17096);
	not 	XG8729 	(g19732,g17096);
	not 	XG8730 	(g19712,g17096);
	not 	XG8731 	(g19687,g17096);
	not 	XG8732 	(g19742,g17096);
	not 	XG8733 	(g19787,g17096);
	not 	XG8734 	(g19743,g17125);
	not 	XG8735 	(g20025,g17271);
	not 	XG8736 	(g19996,g17271);
	not 	XG8737 	(g20533,g17271);
	not 	XG8738 	(g20026,g17271);
	not 	XG8739 	(g19878,g17271);
	not 	XG8740 	(g20040,g17271);
	not 	XG8741 	(I20937,g16967);
	not 	XG8742 	(I20584,g16587);
	not 	XG8743 	(I21210,g17526);
	not 	XG8744 	(g20555,g15480);
	not 	XG8745 	(g21204,g15656);
	not 	XG8746 	(g21205,g15656);
	not 	XG8747 	(g21252,g15656);
	not 	XG8748 	(g20737,g15656);
	not 	XG8749 	(g18880,g15656);
	not 	XG8750 	(g21155,g15656);
	not 	XG8751 	(I19796,g17870);
	not 	XG8752 	(g20625,g15348);
	not 	XG8753 	(g20514,g15348);
	not 	XG8754 	(g20435,g15348);
	not 	XG8755 	(g20538,g15348);
	not 	XG8756 	(g20554,g15348);
	not 	XG8757 	(g20680,g15348);
	not 	XG8758 	(g20650,g15348);
	not 	XG8759 	(g20498,g15348);
	not 	XG8760 	(g20600,g15348);
	not 	XG8761 	(g21461,g15348);
	not 	XG8762 	(g19885,g17249);
	not 	XG8763 	(g20903,g17249);
	not 	XG8764 	(g20004,g17249);
	not 	XG8765 	(g20656,g17249);
	not 	XG8766 	(g20087,g17249);
	not 	XG8767 	(g20579,g17249);
	not 	XG8768 	(g20179,g17249);
	not 	XG8769 	(g19747,g17015);
	not 	XG8770 	(g20247,g17015);
	not 	XG8771 	(g19695,g17015);
	not 	XG8772 	(g20207,g17015);
	not 	XG8773 	(g19776,g17015);
	not 	XG8774 	(g19629,g17015);
	not 	XG8775 	(g19777,g17015);
	not 	XG8776 	(g19718,g17015);
	not 	XG8777 	(g19649,g17015);
	not 	XG8778 	(g19760,g17015);
	not 	XG8779 	(g19682,g17015);
	not 	XG8780 	(g19789,g17015);
	not 	XG8781 	(g19761,g17015);
	not 	XG8782 	(g19852,g17015);
	not 	XG8783 	(g19748,g17015);
	not 	XG8784 	(g20229,g17015);
	not 	XG8785 	(g19696,g17015);
	not 	XG8786 	(g19737,g17015);
	not 	XG8787 	(g20320,g17015);
	not 	XG8788 	(g19872,g17015);
	not 	XG8789 	(g19790,g16971);
	not 	XG8790 	(g20190,g16971);
	not 	XG8791 	(g19698,g16971);
	not 	XG8792 	(g20167,g16971);
	not 	XG8793 	(g20158,g16971);
	not 	XG8794 	(g19650,g16971);
	not 	XG8795 	(g20178,g16971);
	not 	XG8796 	(I21006,g15579);
	not 	XG8797 	(I20913,g16964);
	not 	XG8798 	(I21115,g15714);
	not 	XG8799 	(g20191,g17821);
	not 	XG8800 	(g20541,g17821);
	not 	XG8801 	(g21346,g17821);
	not 	XG8802 	(g21355,g17821);
	not 	XG8803 	(g20379,g17821);
	not 	XG8804 	(g20209,g17821);
	not 	XG8805 	(g21418,g17821);
	not 	XG8806 	(g20523,g17821);
	not 	XG8807 	(g20265,g17821);
	not 	XG8808 	(g20321,g17821);
	not 	XG8809 	(g20231,g17821);
	not 	XG8810 	(g20103,g17433);
	not 	XG8811 	(g20766,g17433);
	not 	XG8812 	(g20005,g17433);
	not 	XG8813 	(g20036,g17433);
	not 	XG8814 	(g20657,g17433);
	not 	XG8815 	(g20697,g17433);
	not 	XG8816 	(g20627,g17433);
	not 	XG8817 	(g20104,g17433);
	not 	XG8818 	(g20090,g17433);
	not 	XG8819 	(g21049,g17433);
	not 	XG8820 	(g20105,g17433);
	not 	XG8821 	(g19960,g17433);
	not 	XG8822 	(g20904,g17433);
	not 	XG8823 	(g20601,g17433);
	not 	XG8824 	(g20066,g17433);
	not 	XG8825 	(g20067,g17328);
	not 	XG8826 	(g20147,g17328);
	not 	XG8827 	(g20106,g17328);
	not 	XG8828 	(g20560,g17328);
	not 	XG8829 	(g20053,g17328);
	not 	XG8830 	(g20037,g17328);
	not 	XG8831 	(g20079,g17328);
	not 	XG8832 	(g20080,g17328);
	not 	XG8833 	(g20129,g17328);
	not 	XG8834 	(g20091,g17328);
	not 	XG8835 	(g20006,g17328);
	not 	XG8836 	(g20130,g17328);
	not 	XG8837 	(g19961,g17328);
	not 	XG8838 	(g20580,g17328);
	not 	XG8839 	(g19912,g17328);
	not 	XG8840 	(g20038,g17328);
	not 	XG8841 	(g20054,g17328);
	not 	XG8842 	(I20529,g16309);
	not 	XG8843 	(g20157,g16886);
	not 	XG8844 	(g20166,g16886);
	not 	XG8845 	(g19697,g16886);
	not 	XG8846 	(g20102,g17533);
	not 	XG8847 	(g20088,g17533);
	not 	XG8848 	(g20089,g17533);
	not 	XG8849 	(g20146,g17533);
	not 	XG8850 	(g20052,g17533);
	not 	XG8851 	(g20064,g17533);
	not 	XG8852 	(g20101,g17533);
	not 	XG8853 	(g20144,g17533);
	not 	XG8854 	(g20159,g17533);
	not 	XG8855 	(g20696,g17533);
	not 	XG8856 	(g20145,g17533);
	not 	XG8857 	(g20128,g17533);
	not 	XG8858 	(g21048,g17533);
	not 	XG8859 	(g20208,g17533);
	not 	XG8860 	(g21295,g17533);
	not 	XG8861 	(g20168,g17533);
	not 	XG8862 	(g20180,g17533);
	not 	XG8863 	(g20671,g15509);
	not 	XG8864 	(g21182,g15509);
	not 	XG8865 	(g18889,g15509);
	not 	XG8866 	(g21249,g15509);
	not 	XG8867 	(g20591,g15509);
	not 	XG8868 	(g21183,g15509);
	not 	XG8869 	(g20507,g15509);
	not 	XG8870 	(g21286,g15509);
	not 	XG8871 	(g20712,g15509);
	not 	XG8872 	(g21456,g15509);
	not 	XG8873 	(g21060,g15509);
	not 	XG8874 	(g21059,g15509);
	not 	XG8875 	(g20529,g15509);
	not 	XG8876 	(g20448,g15509);
	not 	XG8877 	(g18897,g15509);
	not 	XG8878 	(g20779,g15509);
	not 	XG8879 	(g20710,g15509);
	not 	XG8880 	(g20780,g15509);
	not 	XG8881 	(g21184,g15509);
	not 	XG8882 	(g20711,g15509);
	not 	XG8883 	(g20641,g15509);
	not 	XG8884 	(g20530,g15509);
	not 	XG8885 	(g21466,g15509);
	not 	XG8886 	(g20615,g15509);
	not 	XG8887 	(g20568,g15509);
	not 	XG8888 	(g21425,g15509);
	not 	XG8889 	(g21380,g17955);
	not 	XG8890 	(g20562,g17955);
	not 	XG8891 	(g21396,g17955);
	not 	XG8892 	(g20629,g17955);
	not 	XG8893 	(g20701,g17955);
	not 	XG8894 	(g20324,g17955);
	not 	XG8895 	(g20770,g17955);
	not 	XG8896 	(g18828,g17955);
	not 	XG8897 	(g20605,g17955);
	not 	XG8898 	(g20585,g17955);
	not 	XG8899 	(g21178,g17955);
	not 	XG8900 	(g20501,g17955);
	not 	XG8901 	(g20630,g17955);
	not 	XG8902 	(g20267,g17955);
	not 	XG8903 	(g20525,g17955);
	not 	XG8904 	(g20380,g17955);
	not 	XG8905 	(g21406,g17955);
	not 	XG8906 	(g20768,g17955);
	not 	XG8907 	(g20769,g17955);
	not 	XG8908 	(g21608,g17955);
	not 	XG8909 	(g20702,g17955);
	not 	XG8910 	(g20381,g17955);
	not 	XG8911 	(g20606,g17955);
	not 	XG8912 	(g20607,g17955);
	not 	XG8913 	(g20543,g17955);
	not 	XG8914 	(g20909,g17955);
	not 	XG8915 	(I20562,g16525);
	not 	XG8916 	(g19676,g17062);
	not 	XG8917 	(g19659,g17062);
	not 	XG8918 	(g19754,g17062);
	not 	XG8919 	(g19770,g17062);
	not 	XG8920 	(g19799,g17062);
	not 	XG8921 	(g19686,g17062);
	not 	XG8922 	(g20213,g17062);
	not 	XG8923 	(g19730,g17062);
	not 	XG8924 	(g19786,g17062);
	not 	XG8925 	(g19711,g17062);
	not 	XG8926 	(I20895,g16954);
	not 	XG8927 	(g19979,g17226);
	not 	XG8928 	(g19860,g17226);
	not 	XG8929 	(g19980,g17226);
	not 	XG8930 	(g19947,g17226);
	not 	XG8931 	(g20010,g17226);
	not 	XG8932 	(g20510,g17226);
	not 	XG8933 	(g19731,g17093);
	not 	XG8934 	(g19409,g16431);
	not 	XG8935 	(g19763,g16431);
	not 	XG8936 	(g19395,g16431);
	not 	XG8937 	(g19477,g16431);
	not 	XG8938 	(g19386,g16431);
	not 	XG8939 	(g19387,g16431);
	not 	XG8940 	(g19779,g16431);
	not 	XG8941 	(g19396,g16431);
	not 	XG8942 	(g19468,g15938);
	not 	XG8943 	(g19451,g15938);
	not 	XG8944 	(g18883,g15938);
	not 	XG8945 	(g18874,g15938);
	not 	XG8946 	(g21604,g15938);
	not 	XG8947 	(g18944,g15938);
	not 	XG8948 	(g19558,g15938);
	not 	XG8949 	(g18884,g15938);
	not 	XG8950 	(g18975,g15938);
	not 	XG8951 	(g19537,g15938);
	not 	XG8952 	(g19539,g16129);
	not 	XG8953 	(g19577,g16129);
	not 	XG8954 	(g19559,g16129);
	not 	XG8955 	(g19523,g16100);
	not 	XG8956 	(g18946,g16100);
	not 	XG8957 	(g19273,g16100);
	not 	XG8958 	(g19538,g16100);
	not 	XG8959 	(g18976,g16100);
	not 	XG8960 	(g18977,g16100);
	not 	XG8961 	(g18945,g16100);
	not 	XG8962 	(g18929,g16100);
	not 	XG8963 	(g18908,g16100);
	not 	XG8964 	(g19670,g16897);
	not 	XG8965 	(g19612,g16897);
	not 	XG8966 	(g19719,g16897);
	not 	XG8967 	(g20194,g16897);
	not 	XG8968 	(g19652,g16897);
	not 	XG8969 	(g19653,g16897);
	not 	XG8970 	(g19630,g16897);
	not 	XG8971 	(g20182,g16897);
	not 	XG8972 	(g19765,g16897);
	not 	XG8973 	(g20110,g16897);
	not 	XG8974 	(g20210,g16897);
	not 	XG8975 	(g19762,g16326);
	not 	XG8976 	(g19469,g16326);
	not 	XG8977 	(g19385,g16326);
	not 	XG8978 	(g19394,g16326);
	not 	XG8979 	(g19434,g16326);
	not 	XG8980 	(g19421,g16326);
	not 	XG8981 	(g19963,g16326);
	not 	XG8982 	(g19476,g16326);
	not 	XG8983 	(g19368,g16326);
	not 	XG8984 	(g19452,g16326);
	not 	XG8985 	(g19750,g16326);
	not 	XG8986 	(g18885,g15979);
	not 	XG8987 	(g19067,g15979);
	not 	XG8988 	(g18907,g15979);
	not 	XG8989 	(g18988,g15979);
	not 	XG8990 	(g19542,g16349);
	not 	XG8991 	(g19437,g16349);
	not 	XG8992 	(g19493,g16349);
	not 	XG8993 	(g19586,g16349);
	not 	XG8994 	(g19569,g16349);
	not 	XG8995 	(g19543,g16349);
	not 	XG8996 	(g19618,g16349);
	not 	XG8997 	(g19480,g16349);
	not 	XG8998 	(g19526,g16349);
	not 	XG8999 	(g19503,g16349);
	not 	XG9000 	(g19527,g16349);
	not 	XG9001 	(g19481,g16349);
	not 	XG9002 	(g19472,g16349);
	not 	XG9003 	(g19491,g16349);
	not 	XG9004 	(g20009,g16349);
	not 	XG9005 	(g19473,g16349);
	not 	XG9006 	(g19414,g16349);
	not 	XG9007 	(g19570,g16349);
	not 	XG9008 	(g19454,g16349);
	not 	XG9009 	(g20057,g16349);
	not 	XG9010 	(g19494,g16349);
	not 	XG9011 	(g19915,g16349);
	not 	XG9012 	(g19617,g16349);
	not 	XG9013 	(g19544,g16349);
	not 	XG9014 	(g19657,g16349);
	not 	XG9015 	(g19602,g16349);
	not 	XG9016 	(g19528,g16349);
	not 	XG9017 	(g19529,g16349);
	not 	XG9018 	(g19504,g16349);
	not 	XG9019 	(g19603,g16349);
	not 	XG9020 	(g19505,g16349);
	not 	XG9021 	(g19482,g16349);
	not 	XG9022 	(g19634,g16349);
	not 	XG9023 	(g19492,g16349);
	not 	XG9024 	(g19635,g16349);
	not 	XG9025 	(g21050,g17873);
	not 	XG9026 	(g21379,g17873);
	not 	XG9027 	(g20659,g17873);
	not 	XG9028 	(g20700,g17873);
	not 	XG9029 	(g20698,g17873);
	not 	XG9030 	(g20699,g17873);
	not 	XG9031 	(g20767,g17873);
	not 	XG9032 	(g20604,g17873);
	not 	XG9033 	(g21607,g17873);
	not 	XG9034 	(g20500,g17873);
	not 	XG9035 	(g21362,g17873);
	not 	XG9036 	(g20584,g17873);
	not 	XG9037 	(g20441,g17873);
	not 	XG9038 	(g20524,g17873);
	not 	XG9039 	(g20266,g17873);
	not 	XG9040 	(g20561,g17873);
	not 	XG9041 	(g20322,g17873);
	not 	XG9042 	(g20323,g17873);
	not 	XG9043 	(g21395,g17873);
	not 	XG9044 	(g20603,g17873);
	not 	XG9045 	(g20582,g17873);
	not 	XG9046 	(g20233,g17873);
	not 	XG9047 	(g20583,g17873);
	not 	XG9048 	(g20542,g17873);
	not 	XG9049 	(g21560,g17873);
	not 	XG9050 	(g20660,g17873);
	not 	XG9051 	(g19431,g16249);
	not 	XG9052 	(g19360,g16249);
	not 	XG9053 	(g19438,g16249);
	not 	XG9054 	(g19365,g16249);
	not 	XG9055 	(I20216,g15862);
	not 	XG9056 	(g20526,g15171);
	not 	XG9057 	(g20910,g15171);
	not 	XG9058 	(g20661,g15171);
	not 	XG9059 	(g20632,g15171);
	not 	XG9060 	(g20911,g15171);
	not 	XG9061 	(g21051,g15171);
	not 	XG9062 	(g21397,g15171);
	not 	XG9063 	(g20633,g15171);
	not 	XG9064 	(g20563,g15171);
	not 	XG9065 	(g20325,g15171);
	not 	XG9066 	(g18829,g15171);
	not 	XG9067 	(g20771,g15171);
	not 	XG9068 	(g20608,g15171);
	not 	XG9069 	(g20382,g15171);
	not 	XG9070 	(g18875,g15171);
	not 	XG9071 	(g20544,g15171);
	not 	XG9072 	(g20631,g15171);
	not 	XG9073 	(g21247,g15171);
	not 	XG9074 	(g21421,g15171);
	not 	XG9075 	(g20662,g15171);
	not 	XG9076 	(g21407,g15171);
	not 	XG9077 	(g20912,g15171);
	not 	XG9078 	(g20442,g15171);
	not 	XG9079 	(g20586,g15171);
	not 	XG9080 	(g20772,g15171);
	not 	XG9081 	(g20443,g15171);
	not 	XG9082 	(g19905,g15885);
	not 	XG9083 	(g19416,g15885);
	not 	XG9084 	(g19366,g15885);
	not 	XG9085 	(g19950,g15885);
	not 	XG9086 	(g19744,g15885);
	not 	XG9087 	(g19439,g15885);
	not 	XG9088 	(g19865,g15885);
	not 	XG9089 	(g19432,g15885);
	not 	XG9090 	(g19678,g16752);
	not 	XG9091 	(g19498,g16752);
	not 	XG9092 	(g19531,g16816);
	not 	XG9093 	(g19713,g16816);
	not 	XG9094 	(g19733,g16856);
	not 	XG9095 	(g19552,g16856);
	not 	XG9096 	(g20551,g17302);
	not 	XG9097 	(g20059,g17302);
	not 	XG9098 	(g18916,g16053);
	not 	XG9099 	(g18938,g16053);
	not 	XG9100 	(g18904,g16053);
	not 	XG9101 	(g18891,g16053);
	not 	XG9102 	(g18952,g16053);
	not 	XG9103 	(g19517,g16777);
	not 	XG9104 	(g19688,g16777);
	not 	XG9105 	(g20058,g16782);
	not 	XG9106 	(g20096,g16782);
	not 	XG9107 	(g19679,g16782);
	not 	XG9108 	(g19499,g16782);
	not 	XG9109 	(g20153,g16782);
	not 	XG9110 	(g19553,g16782);
	not 	XG9111 	(g20597,g17847);
	not 	XG9112 	(g20240,g17847);
	not 	XG9113 	(g20535,g17847);
	not 	XG9114 	(g20494,g17847);
	not 	XG9115 	(g20432,g17847);
	not 	XG9116 	(g20552,g17847);
	not 	XG9117 	(g21400,g17847);
	not 	XG9118 	(g20574,g17847);
	not 	XG9119 	(g20274,g17847);
	not 	XG9120 	(g20372,g17847);
	not 	XG9121 	(g20495,g17926);
	not 	XG9122 	(I19756,g17812);
	not 	XG9123 	(I21181,g17413);
	not 	XG9124 	(g20978,g15595);
	not 	XG9125 	(g20732,g15595);
	not 	XG9126 	(g20852,g15595);
	not 	XG9127 	(g20622,g15595);
	not 	XG9128 	(g20853,g15595);
	not 	XG9129 	(g21561,g15595);
	not 	XG9130 	(g19373,g16449);
	not 	XG9131 	(g19479,g16449);
	not 	XG9132 	(g19410,g16449);
	not 	XG9133 	(g19443,g16449);
	not 	XG9134 	(g19766,g16449);
	not 	XG9135 	(g20008,g16449);
	not 	XG9136 	(g19435,g16449);
	not 	XG9137 	(g19489,g16449);
	not 	XG9138 	(g19471,g16449);
	not 	XG9139 	(g19780,g16449);
	not 	XG9140 	(g19397,g16449);
	not 	XG9141 	(g19565,g16000);
	not 	XG9142 	(g18978,g16000);
	not 	XG9143 	(g18894,g16000);
	not 	XG9144 	(g19579,g16000);
	not 	XG9145 	(g18895,g16000);
	not 	XG9146 	(g19478,g16000);
	not 	XG9147 	(g18886,g16000);
	not 	XG9148 	(g18989,g16000);
	not 	XG9149 	(g19470,g16000);
	not 	XG9150 	(g18827,g16000);
	not 	XG9151 	(g18931,g16031);
	not 	XG9152 	(g18896,g16031);
	not 	XG9153 	(g19144,g16031);
	not 	XG9154 	(g19068,g16031);
	not 	XG9155 	(g20211,g16931);
	not 	XG9156 	(g19654,g16931);
	not 	XG9157 	(g19739,g16931);
	not 	XG9158 	(g19633,g16931);
	not 	XG9159 	(g20195,g16931);
	not 	XG9160 	(g19683,g16931);
	not 	XG9161 	(g20132,g16931);
	not 	XG9162 	(g20232,g16931);
	not 	XG9163 	(g19783,g16931);
	not 	XG9164 	(g19672,g16931);
	not 	XG9165 	(g19673,g16931);
	not 	XG9166 	(g19781,g16489);
	not 	XG9167 	(g19411,g16489);
	not 	XG9168 	(g19490,g16489);
	not 	XG9169 	(g19794,g16489);
	not 	XG9170 	(g19398,g16489);
	not 	XG9171 	(g19399,g16489);
	not 	XG9172 	(g19429,g16489);
	not 	XG9173 	(g19412,g16489);
	not 	XG9174 	(g18979,g16136);
	not 	XG9175 	(g18980,g16136);
	not 	XG9176 	(g18990,g16136);
	not 	XG9177 	(g18947,g16136);
	not 	XG9178 	(g18991,g16136);
	not 	XG9179 	(g19541,g16136);
	not 	XG9180 	(g19566,g16136);
	not 	XG9181 	(g18932,g16136);
	not 	XG9182 	(g19343,g16136);
	not 	XG9183 	(g19600,g16164);
	not 	XG9184 	(g19580,g16164);
	not 	XG9185 	(g19567,g16164);
	not 	XG9186 	(I21067,g15573);
	not 	XG9187 	(g21428,g15758);
	not 	XG9188 	(g21412,g15758);
	not 	XG9189 	(g18903,g15758);
	not 	XG9190 	(g19415,g15758);
	not 	XG9191 	(g19352,g15758);
	not 	XG9192 	(g21349,g15758);
	not 	XG9193 	(g21305,g15758);
	not 	XG9194 	(g21467,g15758);
	not 	XG9195 	(g21458,g15758);
	not 	XG9196 	(g21337,g15758);
	not 	XG9197 	(g20273,g17128);
	not 	XG9198 	(g20239,g17128);
	not 	XG9199 	(I20690,g15733);
	not 	XG9200 	(g19772,g17183);
	not 	XG9201 	(g20534,g17183);
	not 	XG9202 	(g19208,g17367);
	not 	XG9203 	(g19351,g17367);
	not 	XG9204 	(g21457,g17367);
	not 	XG9205 	(g21427,g17367);
	not 	XG9206 	(g19276,g17367);
	not 	XG9207 	(g21304,g17367);
	not 	XG9208 	(g21383,g17367);
	not 	XG9209 	(g21336,g17367);
	not 	XG9210 	(g18832,g15634);
	not 	XG9211 	(g20679,g15634);
	not 	XG9212 	(g21138,g15634);
	not 	XG9213 	(g21139,g15634);
	not 	XG9214 	(g21189,g15634);
	not 	XG9215 	(g21010,g15634);
	not 	XG9216 	(I19786,g17844);
	not 	XG9217 	(I21199,g17501);
	not 	XG9218 	(g20537,g15345);
	not 	XG9219 	(g20624,g18065);
	not 	XG9220 	(g20497,g18065);
	not 	XG9221 	(g20649,g18065);
	not 	XG9222 	(g20434,g18065);
	not 	XG9223 	(g20576,g18065);
	not 	XG9224 	(g21431,g18065);
	not 	XG9225 	(g20374,g18065);
	not 	XG9226 	(g20599,g18065);
	not 	XG9227 	(g20513,g18065);
	not 	XG9228 	(g20536,g18065);
	not 	XG9229 	(g20706,g18008);
	not 	XG9230 	(g20384,g18008);
	not 	XG9231 	(g20707,g18008);
	not 	XG9232 	(g20527,g18008);
	not 	XG9233 	(g20546,g18008);
	not 	XG9234 	(g20385,g18008);
	not 	XG9235 	(g20776,g18008);
	not 	XG9236 	(g20612,g18008);
	not 	XG9237 	(g21381,g18008);
	not 	XG9238 	(g21409,g18008);
	not 	XG9239 	(g20636,g18008);
	not 	XG9240 	(g21180,g18008);
	not 	XG9241 	(g20588,g18008);
	not 	XG9242 	(g20610,g18008);
	not 	XG9243 	(g18830,g18008);
	not 	XG9244 	(g20774,g18008);
	not 	XG9245 	(g20611,g18008);
	not 	XG9246 	(g20775,g18008);
	not 	XG9247 	(g20504,g18008);
	not 	XG9248 	(g21398,g18008);
	not 	XG9249 	(g21609,g18008);
	not 	XG9250 	(g20326,g18008);
	not 	XG9251 	(g20635,g18008);
	not 	XG9252 	(g20565,g18008);
	not 	XG9253 	(g20268,g18008);
	not 	XG9254 	(g20916,g18008);
	not 	XG9255 	(I20542,g16508);
	not 	XG9256 	(I20846,g16923);
	not 	XG9257 	(g19710,g17059);
	not 	XG9258 	(g20197,g16987);
	not 	XG9259 	(g19685,g16987);
	not 	XG9260 	(g19741,g16987);
	not 	XG9261 	(g19658,g16987);
	not 	XG9262 	(g19785,g16987);
	not 	XG9263 	(g19636,g16987);
	not 	XG9264 	(g19675,g16987);
	not 	XG9265 	(g19709,g16987);
	not 	XG9266 	(g19753,g16987);
	not 	XG9267 	(g19769,g16987);
	not 	XG9268 	(g19964,g17200);
	not 	XG9269 	(g19930,g17200);
	not 	XG9270 	(g19931,g17200);
	not 	XG9271 	(g19902,g17200);
	not 	XG9272 	(g19798,g17200);
	not 	XG9273 	(g20452,g17200);
	not 	XG9274 	(g20917,g15224);
	not 	XG9275 	(g18877,g15224);
	not 	XG9276 	(g20547,g15224);
	not 	XG9277 	(g21248,g15224);
	not 	XG9278 	(g20446,g15224);
	not 	XG9279 	(g20777,g15224);
	not 	XG9280 	(g20613,g15224);
	not 	XG9281 	(g21423,g15224);
	not 	XG9282 	(g20566,g15224);
	not 	XG9283 	(g21410,g15224);
	not 	XG9284 	(g20637,g15224);
	not 	XG9285 	(g20589,g15224);
	not 	XG9286 	(g21055,g15224);
	not 	XG9287 	(g20918,g15224);
	not 	XG9288 	(g20919,g15224);
	not 	XG9289 	(g20528,g15224);
	not 	XG9290 	(g20445,g15224);
	not 	XG9291 	(g18831,g15224);
	not 	XG9292 	(g20386,g15224);
	not 	XG9293 	(g20778,g15224);
	not 	XG9294 	(g21399,g15224);
	not 	XG9295 	(g20327,g15224);
	not 	XG9296 	(g20638,g15224);
	not 	XG9297 	(g20639,g15224);
	not 	XG9298 	(g20666,g15224);
	not 	XG9299 	(g20667,g15224);
	not 	XG9300 	(g20923,g15277);
	not 	XG9301 	(g20450,g15277);
	not 	XG9302 	(g20714,g15277);
	not 	XG9303 	(g20715,g15277);
	not 	XG9304 	(g20451,g15277);
	not 	XG9305 	(g20389,g15277);
	not 	XG9306 	(g20235,g15277);
	not 	XG9307 	(g20329,g15277);
	not 	XG9308 	(g20674,g15277);
	not 	XG9309 	(g20594,g15277);
	not 	XG9310 	(g20570,g15277);
	not 	XG9311 	(g20642,g15277);
	not 	XG9312 	(g20616,g15277);
	not 	XG9313 	(g20617,g15277);
	not 	XG9314 	(g20270,g15277);
	not 	XG9315 	(g20713,g15277);
	not 	XG9316 	(g21426,g15277);
	not 	XG9317 	(g20571,g15277);
	not 	XG9318 	(g20532,g15277);
	not 	XG9319 	(g20549,g15277);
	not 	XG9320 	(g20716,g15277);
	not 	XG9321 	(g20449,g15277);
	not 	XG9322 	(g20672,g15277);
	not 	XG9323 	(g20592,g15277);
	not 	XG9324 	(g20508,g15277);
	not 	XG9325 	(g20509,g15277);
	not 	XG9326 	(g20673,g15277);
	not 	XG9327 	(g21185,g15277);
	not 	XG9328 	(g20593,g15277);
	not 	XG9329 	(g20569,g15277);
	not 	XG9330 	(g20618,g15277);
	not 	XG9331 	(g21068,g15277);
	not 	XG9332 	(g21069,g15277);
	not 	XG9333 	(g20496,g17929);
	not 	XG9334 	(g20623,g17929);
	not 	XG9335 	(g20598,g17929);
	not 	XG9336 	(g20433,g17929);
	not 	XG9337 	(g21414,g17929);
	not 	XG9338 	(g20553,g17929);
	not 	XG9339 	(g20575,g17929);
	not 	XG9340 	(g20275,g17929);
	not 	XG9341 	(g20373,g17929);
	not 	XG9342 	(g20511,g17929);
	not 	XG9343 	(I21189,g17475);
	not 	XG9344 	(I19772,g17818);
	not 	XG9345 	(g20648,g15615);
	not 	XG9346 	(g21123,g15615);
	not 	XG9347 	(g20994,g15615);
	not 	XG9348 	(g20869,g15615);
	not 	XG9349 	(g21610,g15615);
	not 	XG9350 	(g20993,g15615);
	not 	XG9351 	(g20512,g18062);
	not 	XG9352 	(g19952,g15915);
	not 	XG9353 	(g19370,g15915);
	not 	XG9354 	(g19440,g15915);
	not 	XG9355 	(g19755,g15915);
	not 	XG9356 	(g19445,g15915);
	not 	XG9357 	(g19433,g15915);
	not 	XG9358 	(g19998,g15915);
	not 	XG9359 	(g19881,g15915);
	not 	XG9360 	(g19573,g16877);
	not 	XG9361 	(g19745,g16877);
	not 	XG9362 	(g19689,g16795);
	not 	XG9363 	(g19519,g16795);
	not 	XG9364 	(g18917,g16077);
	not 	XG9365 	(g18939,g16077);
	not 	XG9366 	(g18905,g16077);
	not 	XG9367 	(g18983,g16077);
	not 	XG9368 	(g18953,g16077);
	not 	XG9369 	(g19714,g16821);
	not 	XG9370 	(g19532,g16821);
	not 	XG9371 	(g20573,g17384);
	not 	XG9372 	(g20072,g17384);
	not 	XG9373 	(g19734,g16861);
	not 	XG9374 	(g19554,g16861);
	not 	XG9375 	(g20071,g16826);
	not 	XG9376 	(g19520,g16826);
	not 	XG9377 	(g20113,g16826);
	not 	XG9378 	(g20164,g16826);
	not 	XG9379 	(g19690,g16826);
	not 	XG9380 	(g19574,g16826);
	not 	XG9381 	(g21057,g15426);
	not 	XG9382 	(g20590,g15426);
	not 	XG9383 	(g18888,g15426);
	not 	XG9384 	(g20447,g15426);
	not 	XG9385 	(g20506,g15426);
	not 	XG9386 	(g20920,g15426);
	not 	XG9387 	(g21275,g15426);
	not 	XG9388 	(g20921,g15426);
	not 	XG9389 	(g20567,g15426);
	not 	XG9390 	(g21411,g15426);
	not 	XG9391 	(g20668,g15426);
	not 	XG9392 	(g20669,g15426);
	not 	XG9393 	(g21181,g15426);
	not 	XG9394 	(g21058,g15426);
	not 	XG9395 	(g20708,g15426);
	not 	XG9396 	(g20709,g15426);
	not 	XG9397 	(g18878,g15426);
	not 	XG9398 	(g20548,g15426);
	not 	XG9399 	(g20387,g15426);
	not 	XG9400 	(g20505,g15426);
	not 	XG9401 	(g20640,g15426);
	not 	XG9402 	(g20614,g15426);
	not 	XG9403 	(g21455,g15426);
	not 	XG9404 	(g21424,g15426);
	not 	XG9405 	(g20670,g15426);
	not 	XG9406 	(g21056,g15426);
	not 	XG9407 	(I19813,g17952);
	not 	XG9408 	(g20738,g15483);
	not 	XG9409 	(g20515,g15483);
	not 	XG9410 	(g20539,g15483);
	not 	XG9411 	(g20577,g15483);
	not 	XG9412 	(g21511,g15483);
	not 	XG9413 	(g20499,g15483);
	not 	XG9414 	(g20626,g15483);
	not 	XG9415 	(g20681,g15483);
	not 	XG9416 	(g20651,g15483);
	not 	XG9417 	(g20556,g15483);
	not 	XG9418 	(I19661,g17587);
	not 	XG9419 	(g20578,g15563);
	not 	XG9420 	(g21279,g15680);
	not 	XG9421 	(g21268,g15680);
	not 	XG9422 	(g20874,g15680);
	not 	XG9423 	(g18892,g15680);
	not 	XG9424 	(g21221,g15680);
	not 	XG9425 	(g21267,g15680);
	and 	XG9426 	(g20152,g16727,g11545);
	and 	XG9427 	(g20084,g16609,g11591);
	or 	XG9428 	(g23770,g16868,g20188);
	or 	XG9429 	(g22640,g15613,g18951);
	nand 	XG9430 	(g17581,g14669,g5623,g12029,g5607);
	and 	XG9431 	(g24140,g21654,g17663);
	not 	XG9432 	(g17782,I18788);
	or 	XG9433 	(g21895,g15108,g20135);
	or 	XG9434 	(g21894,g15107,g20112);
	nand 	XG9435 	(g16628,g13902,g3618,g11207,g3602);
	or 	XG9436 	(g23217,g16023,g19588);
	nand 	XG9437 	(g21401,g14695,g17712,g14730,g17755);
	nand 	XG9438 	(g17705,g13902,g3661,g13799,g3586);
	nand 	XG9439 	(g17669,g13902,g3632,g11238,g3570);
	and 	XG9440 	(g23436,g20375,g676);
	and 	XG9441 	(g23885,g19513,g4132);
	nand 	XG9442 	(g17650,g14745,g6315,g12101,g6299);
	not 	XG9443 	(I17919,g14609);
	not 	XG9444 	(I17626,g14582);
	not 	XG9445 	(I18304,g14790);
	not 	XG9446 	(g16428,I17668);
	nand 	XG9447 	(g20201,I20469,I20468);
	nand 	XG9448 	(g15781,g14745,g6329,g12173,g6267);
	nand 	XG9449 	(g21415,g14739,g17740,g14771,g17773);
	not 	XG9450 	(g16286,I17615);
	or 	XG9451 	(g24280,g15109,g23292);
	or 	XG9452 	(g21892,g15104,g19788);
	nand 	XG9453 	(g17668,g13877,g3310,g13765,g3235);
	or 	XG9454 	(g22644,g15632,g18981);
	and 	XG9455 	(g23920,g19549,g4135);
	not 	XG9456 	(g16601,I17783);
	or 	XG9457 	(g23298,g16179,g19693);
	and 	XG9458 	(g23348,g21393,g15570);
	nand 	XG9459 	(g15737,g13210,g7903,g13115,g13240);
	nor 	XG9460 	(g20234,g14207,g17140);
	nor 	XG9461 	(g19436,g14233,g17176);
	or 	XG9462 	(g23318,g16192,g19716);
	not 	XG9463 	(g15588,I17166);
	nand 	XG9464 	(g20216,I20488,I20487);
	or 	XG9465 	(g21897,g15111,g20095);
	or 	XG9466 	(g21900,g15114,g20977);
	and 	XG9467 	(g23957,g19589,g4138);
	or 	XG9468 	(g23346,g16204,g19736);
	and 	XG9469 	(g22158,g19609,g13698);
	not 	XG9470 	(I17557,g14510);
	not 	XG9471 	(g17531,I18476);
	or 	XG9472 	(g23358,g16212,g19746);
	not 	XG9473 	(g15566,I17143);
	not 	XG9474 	(g16620,I17808);
	not 	XG9475 	(g17155,I18205);
	not 	XG9476 	(g16307,I17633);
	and 	XG9477 	(g20581,g15571,g10801);
	not 	XG9478 	(I18245,g14676);
	not 	XG9479 	(g17408,I18341);
	and 	XG9480 	(g24142,g21657,g17700);
	and 	XG9481 	(g21464,g10872,g16181);
	not 	XG9482 	(g16285,I17612);
	nand 	XG9483 	(g17634,g13877,g3281,g11217,g3219);
	not 	XG9484 	(I19778,g17781);
	not 	XG9485 	(g17431,I18376);
	and 	XG9486 	(g21558,g13729,g15904);
	and 	XG9487 	(g21404,g13569,g16069);
	or 	XG9488 	(g22662,g15679,g19069);
	not 	XG9489 	(I21722,g19264);
	not 	XG9490 	(g16429,I17671);
	not 	XG9491 	(I18160,g14441);
	not 	XG9492 	(g24999,g23626);
	nand 	XG9493 	(g23324,g20181,g703);
	and 	XG9494 	(g19560,g10893,g1157,g15832);
	and 	XG9495 	(g23856,g19483,g4116);
	nor 	XG9496 	(g16246,g11169,g13551);
	and 	XG9497 	(g19631,g16093,g1484);
	nand 	XG9498 	(g20184,g13896,g16719,g13918,g16770);
	not 	XG9499 	(g15506,I17131);
	not 	XG9500 	(g19446,I19917);
	not 	XG9501 	(I21222,g18091);
	not 	XG9502 	(g21690,g16540);
	not 	XG9503 	(g20060,g16540);
	not 	XG9504 	(I21258,g16540);
	not 	XG9505 	(g19908,g16540);
	not 	XG9506 	(g21662,g16540);
	not 	XG9507 	(g19866,g16540);
	not 	XG9508 	(g19957,g16540);
	not 	XG9509 	(g21666,g16540);
	not 	XG9510 	(g21694,g16540);
	not 	XG9511 	(g21670,g16540);
	not 	XG9512 	(I21230,g16540);
	not 	XG9513 	(I21242,g16540);
	not 	XG9514 	(g19882,g16540);
	not 	XG9515 	(I21250,g16540);
	not 	XG9516 	(g21682,g16540);
	not 	XG9517 	(I21226,g16540);
	not 	XG9518 	(g19954,g16540);
	not 	XG9519 	(I21246,g16540);
	not 	XG9520 	(g20046,g16540);
	not 	XG9521 	(g21674,g16540);
	not 	XG9522 	(g19869,g16540);
	not 	XG9523 	(I21234,g16540);
	not 	XG9524 	(g20073,g16540);
	not 	XG9525 	(g21686,g16540);
	not 	XG9526 	(g21678,g16540);
	not 	XG9527 	(I21238,g16540);
	not 	XG9528 	(I21254,g16540);
	or 	XG9529 	(g21893,g18655,g20094);
	not 	XG9530 	(g17953,I18861);
	and 	XG9531 	(g21420,g13596,g16093);
	not 	XG9532 	(I18414,g14359);
	not 	XG9533 	(g16322,I17650);
	or 	XG9534 	(g21901,g15115,g21251);
	not 	XG9535 	(g17590,I18523);
	not 	XG9536 	(g22359,g19495);
	not 	XG9537 	(g22407,g19455);
	not 	XG9538 	(g22529,g19549);
	not 	XG9539 	(g22496,g19510);
	and 	XG9540 	(g22457,g21288,g7717,g7753);
	and 	XG9541 	(g22369,g20783,g7717,g9354);
	not 	XG9542 	(g23234,g20375);
	and 	XG9543 	(g19540,g15904,g1124);
	not 	XG9544 	(I17395,g12952);
	not 	XG9545 	(g17188,I18224);
	and 	XG9546 	(g22384,g20784,g9285,g9354);
	not 	XG9547 	(g22649,g19063);
	or 	XG9548 	(g22547,g20215,g16855);
	nor 	XG9549 	(g16272,g11189,g13580);
	not 	XG9550 	(g16284,I17609);
	and 	XG9551 	(g24143,g21659,g17694);
	not 	XG9552 	(g16600,I17780);
	or 	XG9553 	(g22331,g17809,g21405);
	or 	XG9554 	(g21899,g15113,g20162);
	not 	XG9555 	(I17879,g14386);
	nand 	XG9556 	(g15748,g13241,g7922,g13130,g13257);
	not 	XG9557 	(I18114,g14509);
	or 	XG9558 	(g23194,g19578,g19564);
	not 	XG9559 	(I17569,g14564);
	not 	XG9560 	(I18138,g14277);
	and 	XG9561 	(g23919,g19546,g4122);
	not 	XG9562 	(g15371,I17114);
	not 	XG9563 	(I21047,g17429);
	or 	XG9564 	(g23319,g16193,g19717);
	not 	XG9565 	(g17248,I18262);
	not 	XG9566 	(g15569,I17148);
	not 	XG9567 	(I19775,g17780);
	not 	XG9568 	(I21058,g17747);
	not 	XG9569 	(I21074,g17766);
	not 	XG9570 	(I20355,g17613);
	not 	XG9571 	(I20388,g17724);
	not 	XG9572 	(I20369,g17690);
	or 	XG9573 	(g21891,g15103,g19948);
	not 	XG9574 	(I18191,g14385);
	or 	XG9575 	(g23345,g16203,g19735);
	or 	XG9576 	(g22625,g18933,g18910);
	not 	XG9577 	(g16577,I17747);
	not 	XG9578 	(g22497,g19513);
	not 	XG9579 	(g22408,g19483);
	not 	XG9580 	(g22527,g19546);
	not 	XG9581 	(g22544,g19589);
	or 	XG9582 	(g22679,g15701,g19145);
	or 	XG9583 	(g23296,g16177,g19691);
	not 	XG9584 	(g15169,I17094);
	not 	XG9585 	(I18086,g13856);
	or 	XG9586 	(g23251,g16098,g19637);
	nor 	XG9587 	(g23204,g16488,g19462,g10685);
	nor 	XG9588 	(g23042,g10685,g19462,g16581);
	or 	XG9589 	(g20522,g16893,g691);
	nand 	XG9590 	(g24787,g23079,g3391);
	not 	XG9591 	(I21042,g15824);
	not 	XG9592 	(I19831,g16533);
	not 	XG9593 	(I21013,g15806);
	not 	XG9594 	(I19843,g16594);
	not 	XG9595 	(I19851,g16615);
	not 	XG9596 	(I19863,g16675);
	not 	XG9597 	(I21029,g15816);
	not 	XG9598 	(I19857,g16640);
	or 	XG9599 	(g22645,g15633,g18982);
	and 	XG9600 	(g19596,g16681,g1094);
	and 	XG9601 	(g24378,g22718,g3106);
	nand 	XG9602 	(g16312,g13574,g13580);
	and 	XG9603 	(g22863,g20388,g9547);
	not 	XG9604 	(g22719,I22024);
	and 	XG9605 	(g24482,g23055,g6875);
	nand 	XG9606 	(g16236,g13058,g13554,g13573);
	or 	XG9607 	(g23276,g16161,g19681);
	nor 	XG9608 	(g19388,g14256,g17181);
	nand 	XG9609 	(g16604,g13877,g3267,g11194,g3251);
	and 	XG9610 	(g19651,g16119,g1111);
	nor 	XG9611 	(g20390,g14257,g17182);
	nor 	XG9612 	(g19430,g14220,g17150);
	or 	XG9613 	(g23261,g16125,g19660);
	and 	XG9614 	(g24649,g23733,g6527);
	and 	XG9615 	(g19610,g16069,g1141);
	or 	XG9616 	(g22653,g15654,g18993);
	and 	XG9617 	(g24014,g19063,g7933);
	nand 	XG9618 	(g22312,g19063,g907);
	and 	XG9619 	(g19383,g13223,g16893);
	nand 	XG9620 	(I20461,I20460,g17515);
	and 	XG9621 	(g24416,g22870,g4939);
	and 	XG9622 	(g25448,g22680,g11202);
	or 	XG9623 	(g23297,g16178,g19692);
	and 	XG9624 	(g23884,g19510,g4119);
	not 	XG9625 	(g24603,g23108);
	nor 	XG9626 	(g19444,g14295,g17192);
	and 	XG9627 	(g23836,g19495,g4129);
	nand 	XG9628 	(g25237,g23711,g6434);
	and 	XG9629 	(g22216,g20000,g13660);
	nand 	XG9630 	(g23047,g20000,g482);
	and 	XG9631 	(g20628,g15789,g1046);
	and 	XG9632 	(g23855,g19455,g4112);
	or 	XG9633 	(g23197,g15966,g19571);
	and 	XG9634 	(g24011,g19524,g7939);
	nand 	XG9635 	(g16291,g13545,g13551);
	nor 	XG9636 	(g19401,g14296,g17193);
	or 	XG9637 	(g23822,g16929,g20218);
	and 	XG9638 	(g22588,g20078,g79);
	or 	XG9639 	(g22530,g20171,g16751);
	nor 	XG9640 	(g24720,g19793,g23051,g1322);
	and 	XG9641 	(g24640,g23733,g6509);
	nand 	XG9642 	(g16225,g13043,g13528,g13544);
	and 	XG9643 	(g24008,g19502,g7909);
	and 	XG9644 	(g22342,g21287,g9285,g9354);
	and 	XG9645 	(g22417,g21186,g9285,g7753);
	and 	XG9646 	(g22472,g21289,g9285,g7753);
	and 	XG9647 	(g24796,g23714,g7097);
	and 	XG9648 	(g22209,g20751,g19907);
	nor 	XG9649 	(g20183,g14222,g17152);
	nor 	XG9650 	(g19400,g14206,g17139);
	or 	XG9651 	(g23720,g16801,g20165);
	nand 	XG9652 	(g15741,g14631,g5320,g14490,g5244);
	or 	XG9653 	(g22901,g15745,g19384);
	and 	XG9654 	(g22432,g21187,g7717,g9354);
	and 	XG9655 	(g22498,g21334,g7717,g7753);
	not 	XG9656 	(g19592,I20035);
	or 	XG9657 	(g23153,g15876,g19521);
	or 	XG9658 	(g23171,g15903,g19536);
	or 	XG9659 	(g23087,g15852,g19487);
	and 	XG9660 	(g24785,g23645,g7051);
	nor 	XG9661 	(g25160,g23659,g5390);
	and 	XG9662 	(g21453,g13625,g16713);
	and 	XG9663 	(g21606,g13763,g15959);
	and 	XG9664 	(g21465,g13663,g16155);
	not 	XG9665 	(I20910,g17197);
	and 	XG9666 	(g22193,g20682,g19880);
	or 	XG9667 	(g23129,g15863,g19500);
	or 	XG9668 	(g23383,g16222,g19756);
	and 	XG9669 	(g24758,g23733,g6523);
	and 	XG9670 	(g22665,g20905,g17174);
	or 	XG9671 	(g23716,g20905,g9194);
	and 	XG9672 	(g24545,g23285,g3333);
	and 	XG9673 	(g24607,g23666,g5817);
	nand 	XG9674 	(g15734,g14631,g5290,g12059,g5228);
	or 	XG9675 	(g22708,g15711,g19266);
	not 	XG9676 	(I22918,g21451);
	and 	XG9677 	(g22298,g21012,g19997);
	and 	XG9678 	(g24687,g23666,g5827);
	or 	XG9679 	(g22751,g15716,g19333);
	not 	XG9680 	(g20230,I20499);
	nor 	XG9681 	(g24766,g23132,g3385);
	and 	XG9682 	(g21452,g13624,g16119);
	and 	XG9683 	(g21419,g13595,g16681);
	nand 	XG9684 	(g17520,g14631,g5276,g12002,g5260);
	and 	XG9685 	(g24820,g23978,g13944);
	nor 	XG9686 	(g24953,g12259,g23978,g10262);
	and 	XG9687 	(g25366,g22406,g7733);
	not 	XG9688 	(I19704,g17653);
	not 	XG9689 	(I19734,g17725);
	not 	XG9690 	(I20569,g16486);
	not 	XG9691 	(I19759,g17767);
	not 	XG9692 	(I20495,g16283);
	not 	XG9693 	(I20447,g16244);
	not 	XG9694 	(I19789,g17793);
	or 	XG9695 	(g22641,g15631,g18974);
	or 	XG9696 	(g23615,g20131,g20109);
	and 	XG9697 	(g22685,g20192,g11891);
	nand 	XG9698 	(g23850,g19462,g12185);
	not 	XG9699 	(g25273,g23978);
	not 	XG9700 	(g18930,g15789);
	or 	XG9701 	(g23374,g13514,g19767);
	and 	XG9702 	(g25285,g13061,g22152);
	or 	XG9703 	(g24580,g13096,g22340);
	and 	XG9704 	(g24731,g23733,g6519);
	not 	XG9705 	(g25109,g23666);
	not 	XG9706 	(g25001,g23666);
	not 	XG9707 	(g25092,g23666);
	not 	XG9708 	(g25016,g23666);
	or 	XG9709 	(g22664,g15694,g19139);
	nor 	XG9710 	(g19453,g14316,g17199);
	nand 	XG9711 	(I16778,g12332,g11292);
	or 	XG9712 	(g23209,g19601,g19585);
	or 	XG9713 	(g22591,g18909,g18893);
	not 	XG9714 	(I20412,g16213);
	not 	XG9715 	(I20399,g16205);
	not 	XG9716 	(I20385,g16194);
	not 	XG9717 	(I20609,g16539);
	not 	XG9718 	(I19799,g17817);
	not 	XG9719 	(I20433,g16234);
	not 	XG9720 	(g22860,g20000);
	nand 	XG9721 	(g15752,g14701,g5983,g12129,g5921);
	nand 	XG9722 	(g15787,g14745,g6358,g14575,g6283);
	not 	XG9723 	(I23149,g19061);
	nand 	XG9724 	(g20214,g13967,g16776,g13993,g16854);
	nor 	XG9725 	(g20149,g14185,g17091);
	nor 	XG9726 	(g19413,g14221,g17151);
	or 	XG9727 	(g23795,g16884,g20203);
	not 	XG9728 	(g23331,g20905);
	and 	XG9729 	(g20658,g15800,g1389);
	not 	XG9730 	(g25047,g23733);
	not 	XG9731 	(g25153,g23733);
	not 	XG9732 	(g25036,g23733);
	not 	XG9733 	(g25133,g23733);
	nand 	XG9734 	(g24809,g23132,g19965);
	nand 	XG9735 	(g21432,g14780,g17761,g14820,g17790);
	nand 	XG9736 	(g15742,g14669,g5637,g12093,g5575);
	nand 	XG9737 	(g15780,g14701,g6012,g14549,g5937);
	nand 	XG9738 	(g17608,g14701,g5969,g12067,g5953);
	or 	XG9739 	(g22318,g17783,g21394);
	nand 	XG9740 	(g15751,g14669,g5666,g14522,g5591);
	not 	XG9741 	(g18948,g15800);
	or 	XG9742 	(g22684,g15703,g19206);
	or 	XG9743 	(g22832,g15722,g19354);
	nand 	XG9744 	(g20198,g13927,g16745,g13958,g16813);
	not 	XG9745 	(g25034,g23695);
	and 	XG9746 	(g24730,g23699,g6177);
	and 	XG9747 	(g24387,g22761,g3457);
	and 	XG9748 	(g19581,g10918,g1500,g15843);
	and 	XG9749 	(g20602,g15580,g10803);
	or 	XG9750 	(g24430,g8234,g23151);
	nand 	XG9751 	(g25216,g23678,g6088);
	and 	XG9752 	(g22307,g21163,g20027);
	and 	XG9753 	(g22208,g20739,g19906);
	not 	XG9754 	(g25072,g23630);
	not 	XG9755 	(g24987,g23630);
	not 	XG9756 	(g25000,g23630);
	not 	XG9757 	(g25090,g23630);
	or 	XG9758 	(g23193,g15937,g19556);
	or 	XG9759 	(g23183,g15911,g19545);
	and 	XG9760 	(g22219,g20887,g19953);
	and 	XG9761 	(g24903,g23889,g128);
	and 	XG9762 	(g23062,g20248,g718);
	or 	XG9763 	(g24557,g19207,g22308);
	and 	XG9764 	(g24790,g23681,g7074);
	and 	XG9765 	(g24659,g23590,g5134);
	and 	XG9766 	(g22299,g21024,g19999);
	not 	XG9767 	(g24604,g23112);
	not 	XG9768 	(g24683,g23112);
	not 	XG9769 	(g24587,g23112);
	not 	XG9770 	(g24667,g23112);
	nand 	XG9771 	(g21462,g14829,g17779,g14871,g17816);
	and 	XG9772 	(g19613,g16713,g1437);
	and 	XG9773 	(g24590,g23413,g6154);
	nand 	XG9774 	(g24776,g23052,g3040);
	nand 	XG9775 	(g16660,g13933,g3969,g11225,g3953);
	nand 	XG9776 	(g17732,g13933,g4012,g13824,g3937);
	or 	XG9777 	(g24398,g21296,g23801);
	and 	XG9778 	(g19671,g16155,g1454);
	and 	XG9779 	(g22937,g20540,g753);
	and 	XG9780 	(g24628,g23666,g5835);
	or 	XG9781 	(g22639,g15612,g18950);
	and 	XG9782 	(g24484,g23208,g16288);
	and 	XG9783 	(g23007,g20248,g681);
	and 	XG9784 	(g24922,g23931,g4831);
	and 	XG9785 	(g24421,g23139,g3835);
	not 	XG9786 	(g24795,g23342);
	or 	XG9787 	(g22648,g15652,g18987);
	or 	XG9788 	(g24390,g21285,g23779);
	nand 	XG9789 	(g17706,g13933,g3983,g11255,g3921);
	or 	XG9790 	(g23275,g16160,g19680);
	or 	XG9791 	(g24565,g19275,g22309);
	nand 	XG9792 	(g15798,g14786,g6704,g14602,g6629);
	nand 	XG9793 	(g24528,g22654,g4098);
	and 	XG9794 	(g25229,g22654,g7636);
	or 	XG9795 	(g22634,g15590,g18934);
	and 	XG9796 	(g24411,g22161,g4584);
	and 	XG9797 	(g24713,g23666,g5831);
	not 	XG9798 	(g24985,g23586);
	or 	XG9799 	(g23262,g16126,g19661);
	nand 	XG9800 	(I20462,I20460,g14187);
	and 	XG9801 	(g21513,g10882,g16196);
	or 	XG9802 	(g24401,g21298,g23811);
	or 	XG9803 	(g24443,g21378,g23917);
	and 	XG9804 	(g19568,g15959,g1467);
	or 	XG9805 	(g22636,g15611,g18943);
	and 	XG9806 	(g24475,g23139,g3831);
	not 	XG9807 	(g24665,g23067);
	not 	XG9808 	(g24586,g23067);
	not 	XG9809 	(g24579,g23067);
	not 	XG9810 	(g24655,g23067);
	and 	XG9811 	(g23009,g14219,g20196);
	and 	XG9812 	(g24670,g23590,g5138);
	and 	XG9813 	(g24582,g23402,g5808);
	nand 	XG9814 	(g17689,g14786,g6661,g12137,g6645);
	nor 	XG9815 	(g23871,g21348,g2811);
	and 	XG9816 	(g24930,g23948,g4826);
	nand 	XG9817 	(g21384,g14663,g17675,g14686,g17734);
	nand 	XG9818 	(g25172,g23560,g5052);
	and 	XG9819 	(g24501,g23182,g14000);
	not 	XG9820 	(g24605,g23139);
	not 	XG9821 	(g24626,g23139);
	not 	XG9822 	(g24711,g23139);
	not 	XG9823 	(g24685,g23139);
	nand 	XG9824 	(g25255,g23659,g20979);
	or 	XG9825 	(g20083,g17058,g2902);
	nand 	XG9826 	(g20076,g16521,g13795);
	not 	XG9827 	(g24437,g22654);
	and 	XG9828 	(g23104,g20248,g661);
	not 	XG9829 	(g24585,g23063);
	not 	XG9830 	(g25035,g23699);
	not 	XG9831 	(g25131,g23699);
	not 	XG9832 	(g25111,g23699);
	not 	XG9833 	(g25017,g23699);
	nand 	XG9834 	(g25186,g23602,g5396);
	and 	XG9835 	(g24415,g22869,g4760);
	or 	XG9836 	(g23750,g16840,g20174);
	and 	XG9837 	(g23050,g20248,g655);
	nand 	XG9838 	(g25233,g23623,g20838);
	and 	XG9839 	(g24608,g23425,g6500);
	nor 	XG9840 	(g24701,g19778,g23024,g979);
	and 	XG9841 	(g22218,g20875,g19951);
	nand 	XG9842 	(g25293,g23726,g21190);
	and 	XG9843 	(g24940,g23971,g5011);
	or 	XG9844 	(g25037,g19911,g23103);
	nand 	XG9845 	(g15788,g14786,g6675,g12211,g6613);
	not 	XG9846 	(g23578,I22725);
	not 	XG9847 	(g23620,I22769);
	and 	XG9848 	(g24395,g22845,g4704);
	and 	XG9849 	(g24403,g22858,g4894);
	not 	XG9850 	(g23954,I23099);
	not 	XG9851 	(g24986,g23590);
	not 	XG9852 	(g25070,g23590);
	not 	XG9853 	(g25055,g23590);
	not 	XG9854 	(g24971,g23590);
	or 	XG9855 	(g19534,g13019,g15650);
	not 	XG9856 	(g25202,g23932);
	or 	XG9857 	(g23255,g16122,g19655);
	not 	XG9858 	(g25174,g23890);
	not 	XG9859 	(g25046,g23729);
	not 	XG9860 	(g25327,g22161);
	or 	XG9861 	(g23317,g16191,g19715);
	nand 	XG9862 	(g22325,g19140,g1252);
	and 	XG9863 	(g22142,g19140,g7957);
	or 	XG9864 	(g24432,g21361,g23900);
	nor 	XG9865 	(g25203,g23756,g6428);
	nor 	XG9866 	(g23835,g21303,g2791);
	not 	XG9867 	(g25239,g23972);
	and 	XG9868 	(g22991,g20248,g645);
	or 	XG9869 	(g22659,g15673,g19062);
	nand 	XG9870 	(g23782,g21062,g2741);
	and 	XG9871 	(g22939,g21062,g9708);
	nor 	XG9872 	(g19070,g11720,g16957);
	nand 	XG9873 	(g25334,g23756,g21253);
	not 	XG9874 	(g22660,g19140);
	and 	XG9875 	(g23023,g20248,g650);
	and 	XG9876 	(g22538,g20248,g14035);
	not 	XG9877 	(g25188,g23909);
	not 	XG9878 	(g24789,g23309);
	or 	XG9879 	(g22652,g15653,g18992);
	not 	XG9880 	(g24778,g23286);
	not 	XG9881 	(g23472,g21062);
	and 	XG9882 	(g23130,g20248,g728);
	not 	XG9883 	(g23512,g20248);
	not 	XG9884 	(g23192,g20248);
	not 	XG9885 	(g23530,g20248);
	not 	XG9886 	(g23614,g20248);
	not 	XG9887 	(g23654,g20248);
	not 	XG9888 	(g23550,g20248);
	not 	XG9889 	(g23496,g20248);
	not 	XG9890 	(g23573,g20248);
	and 	XG9891 	(g24392,g23067,g3115);
	and 	XG9892 	(g24436,g23067,g3125);
	and 	XG9893 	(g24569,g23382,g5115);
	nor 	XG9894 	(g25144,g23623,g5046);
	nor 	XG9895 	(g25189,g23726,g6082);
	and 	XG9896 	(g24488,g23082,g6905);
	not 	XG9897 	(g24625,g23135);
	and 	XG9898 	(g24450,g23067,g3129);
	and 	XG9899 	(g24771,g23605,g7028);
	not 	XG9900 	(g25015,g23662);
	nor 	XG9901 	(g23883,g21067,g2779);
	and 	XG9902 	(g24671,g23630,g5481);
	and 	XG9903 	(g24588,g23590,g5142);
	and 	XG9904 	(g24913,g23908,g4821);
	and 	XG9905 	(g24629,g23699,g6163);
	and 	XG9906 	(g24581,g23590,g5124);
	nor 	XG9907 	(g22190,g18949,g2827);
	and 	XG9908 	(g24686,g23630,g5485);
	nand 	XG9909 	(g24814,g23167,g20011);
	and 	XG9910 	(g24572,g23393,g5462);
	nor 	XG9911 	(g23686,g21066,g2767);
	and 	XG9912 	(g24589,g23630,g5471);
	and 	XG9913 	(g24606,g23630,g5489);
	nand 	XG9914 	(g25268,g23692,g21124);
	and 	XG9915 	(g24639,g23699,g6181);
	and 	XG9916 	(g24409,g23112,g3484);
	and 	XG9917 	(g24714,g23699,g6173);
	and 	XG9918 	(g24556,g23341,g4035);
	and 	XG9919 	(g24757,g23563,g7004);
	and 	XG9920 	(g24422,g22896,g4771);
	nor 	XG9921 	(g24751,g23105,g3034);
	and 	XG9922 	(g24464,g23112,g3480);
	nor 	XG9923 	(g23918,g21382,g2799);
	and 	XG9924 	(g24410,g23139,g3817);
	and 	XG9925 	(g24399,g23067,g3133);
	and 	XG9926 	(g24465,g23139,g3827);
	and 	XG9927 	(g24400,g23112,g3466);
	and 	XG9928 	(g24423,g22897,g4950);
	and 	XG9929 	(g24393,g22844,g3808);
	and 	XG9930 	(g24550,g23308,g3684);
	nor 	XG9931 	(g23955,g18890,g2823);
	nand 	XG9932 	(g24804,g23105,g19916);
	or 	XG9933 	(g24842,g22669,g7804);
	nand 	XG9934 	(g24793,g23124,g3742);
	and 	XG9935 	(g24451,g23112,g3476);
	nand 	XG9936 	(g25200,g23642,g5742);
	and 	XG9937 	(g24495,g23127,g6928);
	and 	XG9938 	(g24402,g22857,g4749);
	and 	XG9939 	(g24427,g22919,g4961);
	not 	XG9940 	(g25218,g23949);
	nor 	XG9941 	(g25175,g23692,g5736);
	nor 	XG9942 	(g24779,g23167,g3736);
	nor 	XG9943 	(g23763,g21276,g2795);
	not 	XG9944 	(g18833,I19661);
	not 	XG9945 	(g19277,I19813);
	not 	XG9946 	(g19074,I19772);
	not 	XG9947 	(g21514,I21189);
	and 	XG9948 	(g22310,g20235,g19662);
	not 	XG9949 	(g20785,I20846);
	not 	XG9950 	(g20330,I20542);
	not 	XG9951 	(g21562,I21199);
	not 	XG9952 	(g19147,I19786);
	not 	XG9953 	(g20596,I20690);
	not 	XG9954 	(g21335,I21067);
	not 	XG9955 	(g21468,I21181);
	not 	XG9956 	(g18997,I19756);
	not 	XG9957 	(g19801,I20216);
	not 	XG9958 	(g20924,I20895);
	not 	XG9959 	(g20391,I20562);
	and 	XG9960 	(g23280,g20146,g19417);
	not 	XG9961 	(g20283,I20529);
	and 	XG9962 	(g23220,g20067,g19417);
	not 	XG9963 	(g21387,I21115);
	not 	XG9964 	(g21037,I20913);
	not 	XG9965 	(g21273,I21006);
	not 	XG9966 	(g19210,I19796);
	not 	XG9967 	(g21611,I21210);
	not 	XG9968 	(g20453,I20584);
	not 	XG9969 	(g21070,I20937);
	not 	XG9970 	(g18562,I19384);
	not 	XG9971 	(I22729,g21308);
	not 	XG9972 	(I22485,g21308);
	not 	XG9973 	(I22665,g21308);
	not 	XG9974 	(I21792,g21308);
	not 	XG9975 	(I21802,g21308);
	not 	XG9976 	(I21757,g21308);
	not 	XG9977 	(g23223,g21308);
	not 	XG9978 	(g23211,g21308);
	not 	XG9979 	(I21815,g21308);
	not 	XG9980 	(g23844,g21308);
	not 	XG9981 	(g23789,g21308);
	not 	XG9982 	(I21776,g21308);
	not 	XG9983 	(g23239,g21308);
	not 	XG9984 	(g23865,g21308);
	not 	XG9985 	(g23816,g21308);
	not 	XG9986 	(g23764,g21308);
	not 	XG9987 	(I22692,g21308);
	not 	XG9988 	(I22539,g19606);
	not 	XG9989 	(I22046,g19330);
	not 	XG9990 	(I22422,g19330);
	not 	XG9991 	(I22499,g21160);
	not 	XG9992 	(I22461,g21225);
	not 	XG9993 	(I21959,g20242);
	not 	XG9994 	(g22646,g19389);
	not 	XG9995 	(I22512,g19389);
	not 	XG9996 	(I22458,g18954);
	not 	XG9997 	(g22136,g20277);
	not 	XG9998 	(I22000,g20277);
	not 	XG9999 	(I22380,g21156);
	not 	XG10000 	(g22667,g21156);
	not 	XG10001 	(I22571,g20097);
	not 	XG10002 	(g23267,g20097);
	not 	XG10003 	(I22028,g20204);
	not 	XG10004 	(I22488,g18984);
	not 	XG10005 	(g22137,g21370);
	not 	XG10006 	(I21969,g21370);
	not 	XG10007 	(g22138,g21370);
	not 	XG10008 	(I22425,g19379);
	not 	XG10009 	(g22682,g19379);
	not 	XG10010 	(I22467,g19662);
	not 	XG10011 	(I22444,g19626);
	not 	XG10012 	(I22525,g19345);
	not 	XG10013 	(I21766,g19620);
	not 	XG10014 	(I21849,g19620);
	not 	XG10015 	(I22400,g19620);
	not 	XG10016 	(I22464,g21222);
	not 	XG10017 	(I22542,g19773);
	not 	XG10018 	(I22366,g19757);
	not 	XG10019 	(I22502,g19376);
	not 	XG10020 	(I22331,g19417);
	not 	XG10021 	(I22419,g19638);
	not 	XG10022 	(I21860,g19638);
	not 	XG10023 	(I21784,g19638);
	or 	XG10024 	(g25575,g24140,g24139);
	or 	XG10025 	(g22585,g21061,g20915);
	not 	XG10026 	(I21477,g18695);
	not 	XG10027 	(I21483,g18726);
	or 	XG10028 	(I23163,g21256,g21193,g21127,g20982);
	not 	XG10029 	(g24024,g21193);
	not 	XG10030 	(g24059,g21193);
	not 	XG10031 	(g24045,g21193);
	not 	XG10032 	(g24052,g21193);
	not 	XG10033 	(g24074,g21193);
	not 	XG10034 	(g24031,g21193);
	not 	XG10035 	(I22619,g21193);
	not 	XG10036 	(g24038,g21193);
	not 	XG10037 	(I21297,g18597);
	nor 	XG10038 	(g24148,g19338,g19268);
	not 	XG10039 	(g24150,g19268);
	not 	XG10040 	(I21734,g19268);
	or 	XG10041 	(g25576,g24142,g24141);
	or 	XG10042 	(g22531,g20922,g20773);
	not 	XG10043 	(I21480,g18696);
	or 	XG10044 	(I26523,g21143,g20998,g20857,g20720);
	not 	XG10045 	(g24115,g20998);
	not 	XG10046 	(I22583,g20998);
	not 	XG10047 	(g24101,g20998);
	not 	XG10048 	(g24093,g20998);
	not 	XG10049 	(g24086,g20998);
	not 	XG10050 	(g24079,g20998);
	not 	XG10051 	(g24108,g20998);
	not 	XG10052 	(g24137,g20998);
	not 	XG10053 	(g24130,g20998);
	not 	XG10054 	(g24126,g19935);
	not 	XG10055 	(g24119,g19935);
	not 	XG10056 	(g24075,g19935);
	not 	XG10057 	(g24112,g19935);
	not 	XG10058 	(g24133,g19935);
	not 	XG10059 	(g24097,g19935);
	not 	XG10060 	(g24090,g19935);
	not 	XG10061 	(g24105,g19935);
	not 	XG10062 	(I22114,g19935);
	not 	XG10063 	(g24067,g21256);
	not 	XG10064 	(g24060,g21256);
	not 	XG10065 	(g24025,g21256);
	not 	XG10066 	(g24032,g21256);
	not 	XG10067 	(I22640,g21256);
	not 	XG10068 	(g24053,g21256);
	not 	XG10069 	(g24046,g21256);
	not 	XG10070 	(g24039,g21256);
	not 	XG10071 	(g24127,g19984);
	not 	XG10072 	(g24120,g19984);
	not 	XG10073 	(g24098,g19984);
	not 	XG10074 	(g24134,g19984);
	not 	XG10075 	(g24106,g19984);
	not 	XG10076 	(g24083,g19984);
	not 	XG10077 	(I22131,g19984);
	not 	XG10078 	(g24113,g19984);
	not 	XG10079 	(g24076,g19984);
	or 	XG10080 	(I23162,g20841,g20014,g19968,g19919);
	not 	XG10081 	(g24019,g19968);
	not 	XG10082 	(g24055,g19968);
	not 	XG10083 	(g24048,g19968);
	not 	XG10084 	(I22128,g19968);
	not 	XG10085 	(g24069,g19968);
	not 	XG10086 	(g24062,g19968);
	not 	XG10087 	(g24034,g19968);
	not 	XG10088 	(g24041,g19968);
	not 	XG10089 	(I21288,g18216);
	not 	XG10090 	(I21291,g18273);
	not 	XG10091 	(I22622,g21209);
	not 	XG10092 	(g24088,g21209);
	not 	XG10093 	(g24095,g21209);
	not 	XG10094 	(g24103,g21209);
	not 	XG10095 	(g24124,g21209);
	not 	XG10096 	(g24081,g21209);
	not 	XG10097 	(g24117,g21209);
	not 	XG10098 	(g24110,g21209);
	not 	XG10099 	(g24131,g21209);
	or 	XG10100 	(g25577,g24144,g24143);
	or 	XG10101 	(g23825,g20781,g20705);
	not 	XG10102 	(g24107,g20857);
	not 	XG10103 	(g24100,g20857);
	not 	XG10104 	(g24092,g20857);
	not 	XG10105 	(I22564,g20857);
	not 	XG10106 	(g24078,g20857);
	not 	XG10107 	(g24129,g20857);
	not 	XG10108 	(g24136,g20857);
	not 	XG10109 	(g24122,g20857);
	not 	XG10110 	(g24085,g20857);
	not 	XG10111 	(g24058,g20982);
	not 	XG10112 	(g24029,g20982);
	not 	XG10113 	(g24036,g20982);
	not 	XG10114 	(g24022,g20982);
	not 	XG10115 	(g24065,g20982);
	not 	XG10116 	(g24043,g20982);
	not 	XG10117 	(I22580,g20982);
	not 	XG10118 	(g24072,g20982);
	not 	XG10119 	(g24077,g20720);
	not 	XG10120 	(g24099,g20720);
	not 	XG10121 	(g24121,g20720);
	not 	XG10122 	(g24135,g20720);
	not 	XG10123 	(g24114,g20720);
	not 	XG10124 	(g24128,g20720);
	not 	XG10125 	(I22547,g20720);
	not 	XG10126 	(g24091,g20720);
	not 	XG10127 	(g24084,g20720);
	not 	XG10128 	(g24149,g19338);
	not 	XG10129 	(I21744,g19338);
	nor 	XG10130 	(g24145,g19422,g19402);
	not 	XG10131 	(g24146,g19422);
	not 	XG10132 	(I21787,g19422);
	not 	XG10133 	(g24044,g21127);
	not 	XG10134 	(g24037,g21127);
	not 	XG10135 	(g24030,g21127);
	not 	XG10136 	(g24023,g21127);
	not 	XG10137 	(I22601,g21127);
	not 	XG10138 	(g24051,g21127);
	not 	XG10139 	(g24073,g21127);
	not 	XG10140 	(g24066,g21127);
	not 	XG10141 	(g24102,g21143);
	not 	XG10142 	(g24094,g21143);
	not 	XG10143 	(g24138,g21143);
	not 	XG10144 	(g24087,g21143);
	not 	XG10145 	(g24080,g21143);
	not 	XG10146 	(g24109,g21143);
	not 	XG10147 	(g24116,g21143);
	not 	XG10148 	(I22604,g21143);
	not 	XG10149 	(g24123,g21143);
	not 	XG10150 	(g24147,g19402);
	not 	XG10151 	(I21769,g19402);
	not 	XG10152 	(g24070,g20014);
	not 	XG10153 	(g24049,g20014);
	not 	XG10154 	(g24042,g20014);
	not 	XG10155 	(I22153,g20014);
	not 	XG10156 	(g24056,g20014);
	not 	XG10157 	(g24027,g20014);
	not 	XG10158 	(g24020,g20014);
	not 	XG10159 	(g24063,g20014);
	not 	XG10160 	(g24071,g20841);
	not 	XG10161 	(I22561,g20841);
	not 	XG10162 	(g24028,g20841);
	not 	XG10163 	(g24064,g20841);
	not 	XG10164 	(g24057,g20841);
	not 	XG10165 	(g24050,g20841);
	not 	XG10166 	(g24021,g20841);
	not 	XG10167 	(g24035,g20841);
	not 	XG10168 	(I21294,g18274);
	not 	XG10169 	(g24061,g19919);
	not 	XG10170 	(g24033,g19919);
	not 	XG10171 	(g24068,g19919);
	not 	XG10172 	(g24026,g19919);
	not 	XG10173 	(I22111,g19919);
	not 	XG10174 	(g24047,g19919);
	not 	XG10175 	(g24040,g19919);
	not 	XG10176 	(g24054,g19919);
	not 	XG10177 	(I21285,g18215);
	not 	XG10178 	(I21300,g18598);
	not 	XG10179 	(I21486,g18727);
	not 	XG10180 	(g24111,g19890);
	not 	XG10181 	(g24089,g19890);
	not 	XG10182 	(g24082,g19890);
	not 	XG10183 	(I22096,g19890);
	not 	XG10184 	(g24118,g19890);
	not 	XG10185 	(g24125,g19890);
	not 	XG10186 	(g24132,g19890);
	not 	XG10187 	(g24096,g19890);
	not 	XG10188 	(g24104,g19890);
	not 	XG10189 	(g16920,I18086);
	not 	XG10190 	(g18911,g15169);
	and 	XG10191 	(g23691,g20993,g14731);
	and 	XG10192 	(g23690,g20978,g14726);
	and 	XG10193 	(g25030,g20432,g23251);
	or 	XG10194 	(g21898,g15112,g20152);
	and 	XG10195 	(g24658,g19732,g22645);
	and 	XG10196 	(g25069,g20535,g23296);
	and 	XG10197 	(g24710,g19771,g22679);
	and 	XG10198 	(g24664,g19741,g22652);
	and 	XG10199 	(g25058,g20513,g23276);
	not 	XG10200 	(g21329,g16577);
	and 	XG10201 	(g23606,g20679,g16927);
	and 	XG10202 	(g24618,g19672,g22625);
	and 	XG10203 	(g24748,g22457,g17656);
	and 	XG10204 	(g25108,g20576,g23345);
	not 	XG10205 	(g17141,I18191);
	and 	XG10206 	(g23658,g20852,g14687);
	and 	XG10207 	(g25041,g20494,g23261);
	and 	XG10208 	(g24669,g19742,g22653);
	and 	XG10209 	(g24721,g22369,g17488);
	and 	XG10210 	(g25559,g22649,g13004);
	nand 	XG10211 	(g22687,g7870,g19560);
	nand 	XG10212 	(g22642,g19560,g7870);
	nand 	XG10213 	(g22833,g10666,g19560,g1193);
	nor 	XG10214 	(g22400,g15718,g19345);
	nand 	XG10215 	(g25470,g8365,g2051,g22457);
	and 	XG10216 	(g25449,g22496,g6946);
	and 	XG10217 	(g25367,g22407,g6946);
	not 	XG10218 	(g20100,I20369);
	not 	XG10219 	(g20127,I20388);
	not 	XG10220 	(g20086,I20355);
	not 	XG10221 	(g21340,I21074);
	not 	XG10222 	(g21326,I21058);
	not 	XG10223 	(g19127,I19775);
	not 	XG10224 	(g20041,g15569);
	and 	XG10225 	(g23187,g20010,g13989);
	and 	XG10226 	(g25077,g20536,g23297);
	and 	XG10227 	(g23755,g21204,g14821);
	and 	XG10228 	(g22157,g18892,g14608);
	not 	XG10229 	(g21434,g17248);
	and 	XG10230 	(g24703,g22369,g17592);
	and 	XG10231 	(g23724,g21123,g14767);
	nor 	XG10232 	(g22450,g15724,g19345);
	and 	XG10233 	(g25095,g20556,g23319);
	and 	XG10234 	(g24499,g19394,g22217);
	and 	XG10235 	(g24967,g20213,g23197);
	and 	XG10236 	(g23799,g21279,g14911);
	not 	XG10237 	(g21300,I21047);
	and 	XG10238 	(g23389,g19757,g9072);
	not 	XG10239 	(g20028,g15371);
	and 	XG10240 	(g22899,g19695,g19486);
	and 	XG10241 	(g24723,g22384,g17490);
	and 	XG10242 	(g22622,g19469,g19336);
	not 	XG10243 	(g17010,I18138);
	and 	XG10244 	(g24763,g22457,g17569);
	nand 	XG10245 	(g25389,g12082,g22457);
	nand 	XG10246 	(g25492,g22457,g12479);
	not 	XG10247 	(g16228,I17569);
	and 	XG10248 	(g23372,g20194,g16448);
	and 	XG10249 	(g24962,g20210,g23194);
	and 	XG10250 	(g25551,g21511,g23822);
	and 	XG10251 	(g22831,g19629,g19441);
	and 	XG10252 	(g24673,g19748,g22659);
	not 	XG10253 	(g16960,I18114);
	or 	XG10254 	(g21896,g15110,g20084);
	not 	XG10255 	(I20130,g15748);
	nand 	XG10256 	(g25385,g8241,g1783,g22369);
	not 	XG10257 	(g16677,I17879);
	nor 	XG10258 	(g25005,g23324,g6811);
	nor 	XG10259 	(g25022,g23324,g714);
	and 	XG10260 	(g24532,g19478,g22331);
	not 	XG10261 	(g21299,g16600);
	and 	XG10262 	(g23646,g20737,g16959);
	not 	XG10263 	(I21100,g16284);
	and 	XG10264 	(g24004,g21225,g37);
	nand 	XG10265 	(g25309,g12021,g22384);
	nand 	XG10266 	(g25432,g22384,g12374);
	and 	XG10267 	(g25955,g19580,g24720);
	and 	XG10268 	(g24559,g19567,g22993);
	and 	XG10269 	(g22990,g19760,g19555);
	and 	XG10270 	(g23497,g20569,g20169);
	not 	XG10271 	(g24980,g22384);
	not 	XG10272 	(g25100,g22384);
	not 	XG10273 	(g25101,g22384);
	not 	XG10274 	(g25119,g22384);
	not 	XG10275 	(g24993,g22384);
	not 	XG10276 	(g19666,g17188);
	nand 	XG10277 	(I22944,g19620,g9492);
	not 	XG10278 	(g15932,I17395);
	and 	XG10279 	(g25526,g21400,g23720);
	and 	XG10280 	(g25916,g19434,g24432);
	nor 	XG10281 	(g24959,g23324,g8858);
	nor 	XG10282 	(g24976,g23324,g671);
	and 	XG10283 	(g24803,g20005,g22901);
	not 	XG10284 	(g24979,g22369);
	not 	XG10285 	(g25116,g22369);
	not 	XG10286 	(g24991,g22369);
	not 	XG10287 	(g25098,g22369);
	not 	XG10288 	(g25099,g22369);
	and 	XG10289 	(g23533,g13015,g19436);
	not 	XG10290 	(g25136,g22457);
	not 	XG10291 	(g25007,g22457);
	not 	XG10292 	(g25135,g22457);
	not 	XG10293 	(g25154,g22457);
	not 	XG10294 	(g25023,g22457);
	and 	XG10295 	(g22589,g19451,g19267);
	and 	XG10296 	(g25089,g20553,g23317);
	and 	XG10297 	(g23484,g20541,g20160);
	and 	XG10298 	(g22623,g19470,g19337);
	and 	XG10299 	(g25466,g21346,g23574);
	and 	XG10300 	(g24931,g20178,g23153);
	and 	XG10301 	(g24941,g20190,g23171);
	or 	XG10302 	(g24517,g18906,g22158);
	and 	XG10303 	(g24915,g20158,g23087);
	not 	XG10304 	(I19707,g17590);
	and 	XG10305 	(g23498,g12998,g20234);
	and 	XG10306 	(g22329,g20329,g11940);
	and 	XG10307 	(g23131,g19930,g13919);
	not 	XG10308 	(g21352,g16322);
	not 	XG10309 	(g17487,I18414);
	and 	XG10310 	(g23998,g10971,g19631);
	and 	XG10311 	(g22624,g19471,g19344);
	not 	XG10312 	(g19644,g17953);
	and 	XG10313 	(g24923,g20167,g23129);
	and 	XG10314 	(g23873,g10815,g21222);
	and 	XG10315 	(g23857,g7908,g19626);
	and 	XG10316 	(g23872,g4157,g19389);
	and 	XG10317 	(g25152,g20626,g23383);
	nand 	XG10318 	(g22864,g21156,g7780);
	not 	XG10319 	(g21693,I21254);
	not 	XG10320 	(g21677,I21238);
	not 	XG10321 	(g23203,g20073);
	not 	XG10322 	(g21673,I21234);
	not 	XG10323 	(g23020,g19869);
	not 	XG10324 	(g23170,g20046);
	not 	XG10325 	(g21685,I21246);
	not 	XG10326 	(g23084,g19954);
	not 	XG10327 	(g21665,I21226);
	not 	XG10328 	(g21689,I21250);
	not 	XG10329 	(g23041,g19882);
	not 	XG10330 	(g21681,I21242);
	not 	XG10331 	(g21669,I21230);
	not 	XG10332 	(g23085,g19957);
	not 	XG10333 	(g23019,g19866);
	not 	XG10334 	(g23060,g19908);
	not 	XG10335 	(g21697,I21258);
	not 	XG10336 	(g23189,g20060);
	not 	XG10337 	(g21661,I21222);
	not 	XG10338 	(I22289,g19446);
	not 	XG10339 	(I22286,g19446);
	not 	XG10340 	(g21269,g15506);
	and 	XG10341 	(g23725,g21138,g14772);
	and 	XG10342 	(g26783,g21048,g25037);
	and 	XG10343 	(g24553,g19539,g22983);
	and 	XG10344 	(g25949,g19559,g24701);
	and 	XG10345 	(g23775,g21267,g14872);
	and 	XG10346 	(g23901,g7963,g19606);
	and 	XG10347 	(g23837,g10804,g21160);
	and 	XG10348 	(g23921,g4146,g19379);
	and 	XG10349 	(g23471,g20523,g20148);
	and 	XG10350 	(g23056,g19860,g16052);
	not 	XG10351 	(g17088,I18160);
	and 	XG10352 	(g24743,g19789,g22708);
	and 	XG10353 	(g25530,g21414,g23750);
	and 	XG10354 	(g24761,g19852,g22751);
	not 	XG10355 	(g19694,g16429);
	not 	XG10356 	(g22139,I21722);
	and 	XG10357 	(g24503,g19409,g22225);
	and 	XG10358 	(g22489,g19386,g12954);
	and 	XG10359 	(g22848,g19649,g19449);
	and 	XG10360 	(g22686,g19577,g19335);
	and 	XG10361 	(g23564,g20648,g16882);
	and 	XG10362 	(g23572,g20656,g20230);
	and 	XG10363 	(g24682,g19754,g22662);
	and 	XG10364 	(g22590,g19452,g19274);
	not 	XG10365 	(I19719,g17431);
	and 	XG10366 	(g24012,g21561,g14496);
	not 	XG10367 	(g19128,I19778);
	and 	XG10368 	(g23396,g20229,g20051);
	and 	XG10369 	(g23754,g21189,g14816);
	and 	XG10370 	(g22982,g19747,g19535);
	and 	XG10371 	(g23025,g19798,g16021);
	and 	XG10372 	(g24650,g19718,g22641);
	nand 	XG10373 	(g20133,g14569,g17597,g17634,g17668);
	and 	XG10374 	(g23439,g20452,g13771);
	and 	XG10375 	(g25491,g21355,g23615);
	not 	XG10376 	(g21369,g16285);
	and 	XG10377 	(g23404,g20247,g20063);
	nand 	XG10378 	(I21976,g19620,g7680);
	not 	XG10379 	(I19927,g17408);
	not 	XG10380 	(g17221,I18245);
	or 	XG10381 	(g23989,g17179,g20581);
	and 	XG10382 	(g23008,g19783,g1570);
	and 	XG10383 	(g22862,g19673,g1570);
	not 	XG10384 	(g21358,g16307);
	and 	XG10385 	(g23451,g20510,g13805);
	nand 	XG10386 	(I22972,g19638,g9657);
	not 	XG10387 	(I20781,g17155);
	and 	XG10388 	(g25122,g20592,g23374);
	and 	XG10389 	(g24643,g19696,g22636);
	and 	XG10390 	(g24698,g19761,g22664);
	and 	XG10391 	(g25923,g19443,g24443);
	and 	XG10392 	(g23201,g20040,g14027);
	not 	XG10393 	(g21291,g16620);
	not 	XG10394 	(g18898,g15566);
	nand 	XG10395 	(g23357,g11231,g20201);
	and 	XG10396 	(g25130,g20600,g23358);
	and 	XG10397 	(g25042,g20496,g23262);
	not 	XG10398 	(g21228,g17531);
	and 	XG10399 	(g23387,g20211,g16506);
	and 	XG10400 	(g24977,g20232,g23209);
	and 	XG10401 	(g23373,g20195,g13699);
	and 	XG10402 	(g24600,g19652,g22591);
	not 	XG10403 	(g16216,I17557);
	and 	XG10404 	(g22834,g19630,g102);
	and 	XG10405 	(g24634,g19685,g22634);
	and 	XG10406 	(g23188,g20025,g13994);
	and 	XG10407 	(g22849,g19653,g1227);
	and 	XG10408 	(g22992,g19765,g1227);
	and 	XG10409 	(g25181,g20696,g23405);
	and 	XG10410 	(g25113,g20577,g23346);
	and 	XG10411 	(g22710,g19600,g19358);
	and 	XG10412 	(g24504,g19410,g22226);
	and 	XG10413 	(g26153,g19780,g24565);
	and 	XG10414 	(g23006,g19776,g19575);
	nand 	XG10415 	(g20271,g16628,g16657,g14054,g16925);
	and 	XG10416 	(g25057,g20511,g23275);
	and 	XG10417 	(g23474,g20533,g13830);
	not 	XG10418 	(g21463,g15588);
	and 	XG10419 	(g25543,g21461,g23795);
	and 	XG10420 	(g25900,g19368,g24390);
	and 	XG10421 	(g24660,g19737,g22648);
	nand 	XG10422 	(g20150,g14590,g17635,g17669,g17705);
	and 	XG10423 	(g25094,g20554,g23318);
	not 	XG10424 	(I20116,g15737);
	or 	XG10425 	(g25261,g20193,g23348);
	and 	XG10426 	(g25078,g20538,g23298);
	not 	XG10427 	(g21280,g16601);
	and 	XG10428 	(g23774,g21252,g14867);
	and 	XG10429 	(g24657,g19730,g22644);
	and 	XG10430 	(g23386,g20207,g20034);
	and 	XG10431 	(g23415,g20320,g20077);
	and 	XG10432 	(g23165,g19964,g13954);
	and 	XG10433 	(g24645,g19709,g22639);
	and 	XG10434 	(g22515,g19395,g12981);
	not 	XG10435 	(g21281,g16286);
	and 	XG10436 	(g23397,g20239,g11154);
	and 	XG10437 	(g23407,g20273,g9295);
	nand 	XG10438 	(I21992,g19638,g7670);
	and 	XG10439 	(g23682,g20874,g16970);
	and 	XG10440 	(g25902,g19373,g24398);
	and 	XG10441 	(g22149,g18880,g14581);
	and 	XG10442 	(g22165,g18903,g15594);
	and 	XG10443 	(g22752,g19612,g15792);
	and 	XG10444 	(g22637,g19489,g19363);
	and 	XG10445 	(g22835,g19633,g15803);
	and 	XG10446 	(g22633,g19479,g19359);
	nand 	XG10447 	(g21459,g17581,g17605,g14854,g17814);
	not 	XG10448 	(g21343,g16428);
	and 	XG10449 	(g22851,g19654,g496);
	not 	XG10450 	(g17325,I18304);
	and 	XG10451 	(g23540,g20622,g16866);
	and 	XG10452 	(g26122,g19762,g24557);
	not 	XG10453 	(g16300,I17626);
	and 	XG10454 	(g22316,g20270,g2837);
	not 	XG10455 	(g16709,I17919);
	and 	XG10456 	(g24945,g20197,g23183);
	and 	XG10457 	(g24016,g21610,g14528);
	and 	XG10458 	(g24961,g20209,g23193);
	not 	XG10459 	(g24839,g23436);
	and 	XG10460 	(g22145,g18832,g14555);
	and 	XG10461 	(g22632,g19476,g19356);
	and 	XG10462 	(g22900,g19697,g17137);
	and 	XG10463 	(g24523,g19468,g22318);
	and 	XG10464 	(g23349,g20182,g13662);
	and 	XG10465 	(g24983,g20238,g23217);
	not 	XG10466 	(I20951,g17782);
	and 	XG10467 	(g24507,g19429,g22304);
	nor 	XG10468 	(g22929,g12970,g19773);
	and 	XG10469 	(g22518,g19398,g12982);
	and 	XG10470 	(g22525,g19411,g13006);
	and 	XG10471 	(g23991,g21428,g19209);
	and 	XG10472 	(g23166,g19979,g13959);
	and 	XG10473 	(g24646,g19711,g22640);
	and 	XG10474 	(g23416,g20321,g20082);
	and 	XG10475 	(g25536,g21431,g23770);
	and 	XG10476 	(g24773,g19872,g22832);
	and 	XG10477 	(g24717,g19777,g22684);
	and 	XG10478 	(g23083,g19878,g16076);
	nand 	XG10479 	(g21429,g17520,g17578,g14803,g17788);
	and 	XG10480 	(g25978,g25001,g9391);
	nand 	XG10481 	(g21356,g13118,g15743,g15752,g15780);
	and 	XG10482 	(g24704,g22384,g17593);
	and 	XG10483 	(g24467,g23047,g13761);
	nand 	XG10484 	(g21364,g13131,g15753,g15781,g15787);
	nand 	XG10485 	(g20236,g16604,g16625,g14014,g16875);
	nand 	XG10486 	(g25341,g12047,g22417);
	nor 	XG10487 	(g25004,g23324,g676);
	nor 	XG10488 	(g24990,g23324,g8898);
	nand 	XG10489 	(g21555,g17650,g17686,g14946,g17846);
	or 	XG10490 	(g25941,g22219,g24416);
	and 	XG10491 	(g25815,g24603,g8155);
	not 	XG10492 	(g26083,g24809);
	nand 	XG10493 	(g25400,g12086,g22472);
	nand 	XG10494 	(g21338,g13097,g15728,g15734,g15741);
	nand 	XG10495 	(g25429,g8302,g1917,g22417);
	and 	XG10496 	(g24775,g22498,g17594);
	nand 	XG10497 	(g25498,g8418,g2610,g22498);
	and 	XG10498 	(g25988,g25016,g9510);
	nand 	XG10499 	(g23379,g11248,g20216);
	and 	XG10500 	(g24764,g22472,g17570);
	and 	XG10501 	(g25522,g22544,g6888);
	and 	XG10502 	(g25450,g22497,g6888);
	and 	XG10503 	(g25503,g22529,g6888);
	and 	XG10504 	(g25323,g22359,g6888);
	or 	XG10505 	(g22447,g12761,g21464);
	nand 	XG10506 	(g25435,g8316,g2342,g22432);
	and 	XG10507 	(g24749,g22432,g17511);
	and 	XG10508 	(g25050,g22312,g13056);
	nor 	XG10509 	(g24439,g22312,g7400);
	not 	XG10510 	(g24005,I23149);
	nand 	XG10511 	(I20221,g11170,g16272);
	not 	XG10512 	(g20175,I20433);
	not 	XG10513 	(g19263,I19799);
	not 	XG10514 	(g20516,I20609);
	not 	XG10515 	(g20114,I20385);
	not 	XG10516 	(g20136,I20399);
	not 	XG10517 	(g20154,I20412);
	nand 	XG10518 	(I16780,I16778,g12332);
	and 	XG10519 	(g20069,g8955,g9011,g9051,g16312);
	nand 	XG10520 	(I16779,I16778,g11292);
	nand 	XG10521 	(g25473,g22432,g12437);
	nand 	XG10522 	(g25349,g12051,g22432);
	nand 	XG10523 	(g20200,I20462,I20461);
	and 	XG10524 	(g24724,g22432,g17624);
	and 	XG10525 	(g21559,g10897,g16236);
	nand 	XG10526 	(I20187,g1333,g16272);
	or 	XG10527 	(g25789,g14543,g25285);
	and 	XG10528 	(g21512,g10881,g16225);
	nand 	XG10529 	(I20165,g990,g16246);
	not 	XG10530 	(g24791,g23850);
	and 	XG10531 	(g25975,g24999,g9434);
	not 	XG10532 	(g19200,I19789);
	not 	XG10533 	(g20189,I20447);
	not 	XG10534 	(g20219,I20495);
	not 	XG10535 	(g19050,I19759);
	not 	XG10536 	(g20436,I20569);
	not 	XG10537 	(g18957,I19734);
	not 	XG10538 	(g18918,I19704);
	or 	XG10539 	(g25834,g23854,g25366);
	nand 	XG10540 	(g25426,g22369,g12371);
	nand 	XG10541 	(g25300,g12018,g22369);
	not 	XG10542 	(g26340,g24953);
	nand 	XG10543 	(g25439,g12122,g22498);
	and 	XG10544 	(g24001,g10951,g19651);
	and 	XG10545 	(g23996,g10951,g19596);
	and 	XG10546 	(g23990,g10951,g19610);
	and 	XG10547 	(g24015,g10951,g19540);
	nor 	XG10548 	(g26183,g24766,g23079);
	nand 	XG10549 	(I20203,g11147,g16246);
	nand 	XG10550 	(g25514,g22498,g12540);
	nand 	XG10551 	(g26685,g25160,g9264);
	not 	XG10552 	(g23777,I22918);
	and 	XG10553 	(g20056,g8903,g8954,g9007,g16291);
	nand 	XG10554 	(g25467,g22417,g12432);
	not 	XG10555 	(g24960,g23716);
	or 	XG10556 	(g25929,g22193,g24395);
	and 	XG10557 	(g24722,g22417,g17618);
	or 	XG10558 	(g25936,g22209,g24403);
	nand 	XG10559 	(g25476,g8373,g2476,g22472);
	not 	XG10560 	(g21036,I20910);
	nand 	XG10561 	(g25275,g11991,g22342);
	and 	XG10562 	(g24702,g22342,g17464);
	and 	XG10563 	(g23581,g11900,g20183);
	and 	XG10564 	(g23554,g13024,g20390);
	nand 	XG10565 	(g25396,g8259,g2208,g22384);
	and 	XG10566 	(g24765,g22498,g17699);
	not 	XG10567 	(g25039,g22498);
	not 	XG10568 	(g25156,g22498);
	not 	XG10569 	(g25157,g22498);
	not 	XG10570 	(g25025,g22498);
	not 	XG10571 	(g25170,g22498);
	and 	XG10572 	(g23532,g11852,g19400);
	and 	XG10573 	(g23513,g13007,g19430);
	and 	XG10574 	(g23618,g11917,g19388);
	and 	XG10575 	(g23577,g13033,g19444);
	and 	XG10576 	(g23657,g11941,g19401);
	not 	XG10577 	(g25137,g22432);
	not 	XG10578 	(g25120,g22432);
	not 	XG10579 	(g25121,g22432);
	not 	XG10580 	(g24994,g22432);
	not 	XG10581 	(g25008,g22432);
	or 	XG10582 	(g22872,g19383,g19372);
	and 	XG10583 	(g24750,g22472,g17662);
	not 	XG10584 	(g25024,g22472);
	not 	XG10585 	(g25138,g22472);
	not 	XG10586 	(g25139,g22472);
	not 	XG10587 	(g25009,g22472);
	not 	XG10588 	(g25155,g22472);
	not 	XG10589 	(g25006,g22417);
	not 	XG10590 	(g25117,g22417);
	not 	XG10591 	(g25134,g22417);
	not 	XG10592 	(g25118,g22417);
	not 	XG10593 	(g24992,g22417);
	not 	XG10594 	(g24978,g22342);
	not 	XG10595 	(g24963,g22342);
	not 	XG10596 	(g25082,g22342);
	not 	XG10597 	(g25097,g22342);
	not 	XG10598 	(g25081,g22342);
	or 	XG10599 	(g24496,g21557,g24008);
	or 	XG10600 	(g24500,g21605,g24011);
	or 	XG10601 	(g24746,g19461,g22588);
	not 	XG10602 	(g24699,g23047);
	not 	XG10603 	(I25534,g25448);
	and 	XG10604 	(g25502,g22527,g6946);
	and 	XG10605 	(g25368,g22408,g6946);
	not 	XG10606 	(g25564,g22312);
	or 	XG10607 	(g24896,g19684,g22863);
	not 	XG10608 	(g19371,I19857);
	not 	XG10609 	(g21290,I21029);
	not 	XG10610 	(g19375,I19863);
	not 	XG10611 	(g19367,I19851);
	not 	XG10612 	(g19361,I19843);
	not 	XG10613 	(g21278,I21013);
	not 	XG10614 	(g19353,I19831);
	not 	XG10615 	(g21297,I21042);
	nand 	XG10616 	(g23428,g20522,g13945);
	not 	XG10617 	(g24732,g23042);
	not 	XG10618 	(g24825,g23204);
	not 	XG10619 	(I23711,g23192);
	nand 	XG10620 	(g26235,g24766,g8016);
	and 	XG10621 	(g26078,g25055,g5128);
	and 	XG10622 	(g26085,g25070,g11906);
	and 	XG10623 	(g25881,g24685,g3821);
	and 	XG10624 	(g25884,g24711,g11153);
	nand 	XG10625 	(g25337,g8187,g1648,g22342);
	and 	XG10626 	(g25872,g24655,g3119);
	and 	XG10627 	(g25874,g24665,g11118);
	nand 	XG10628 	(g25495,g22472,g12483);
	and 	XG10629 	(g26077,g25233,g9607);
	and 	XG10630 	(g26120,g25293,g9809);
	and 	XG10631 	(g26097,g25092,g5821);
	and 	XG10632 	(g26119,g25109,g11944);
	and 	XG10633 	(g26050,g25047,g9630);
	and 	XG10634 	(g24573,g23716,g17198);
	and 	XG10635 	(g25967,g24986,g9373);
	nand 	XG10636 	(g22650,g19581,g7888);
	nand 	XG10637 	(g22711,g7888,g19581);
	nand 	XG10638 	(g22850,g10699,g19581,g1536);
	nand 	XG10639 	(g26782,g25203,g9467);
	and 	XG10640 	(g24406,g22860,g13623);
	and 	XG10641 	(g23531,g18930,g10760);
	and 	XG10642 	(g26049,g25046,g9621);
	not 	XG10643 	(g26608,g25334);
	not 	XG10644 	(g25083,g23782);
	and 	XG10645 	(g24675,g22342,g17568);
	nand 	XG10646 	(g25382,g22342,g12333);
	or 	XG10647 	(g22490,g12795,g21513);
	nor 	XG10648 	(g25407,g14645,g23871);
	nor 	XG10649 	(g25321,g14645,g23835);
	and 	XG10650 	(g25976,g25000,g9443);
	and 	XG10651 	(g26021,g25035,g9568);
	or 	XG10652 	(g24935,g19749,g22937);
	and 	XG10653 	(g24747,g22417,g17510);
	and 	XG10654 	(g25816,g24604,g8164);
	nor 	XG10655 	(g26715,g25203,g23711);
	and 	XG10656 	(g25962,g24971,g9258);
	not 	XG10657 	(g24357,g22325);
	and 	XG10658 	(g23619,g13045,g19453);
	and 	XG10659 	(g23553,g11875,g19413);
	nor 	XG10660 	(g24875,g11083,g23850,g8725);
	and 	XG10661 	(g24498,g23850,g14036);
	and 	XG10662 	(g26087,g25072,g5475);
	and 	XG10663 	(g26095,g25090,g11923);
	or 	XG10664 	(g24813,g19594,g22685);
	and 	XG10665 	(g25938,g24953,g8997);
	nand 	XG10666 	(g26382,g12323,g24953,g577);
	and 	XG10667 	(g23514,g11829,g20149);
	or 	XG10668 	(g25942,g22298,g24422);
	nor 	XG10669 	(g26645,g25160,g23602);
	and 	XG10670 	(g26086,g25255,g9672);
	and 	XG10671 	(g24002,g10971,g19613);
	and 	XG10672 	(g22143,g10971,g19568);
	and 	XG10673 	(g24009,g10971,g19671);
	nand 	XG10674 	(g21386,g13139,g15782,g15788,g15798);
	not 	XG10675 	(I24400,g23954);
	and 	XG10676 	(g26147,g25133,g6513);
	and 	XG10677 	(g26165,g25153,g11980);
	not 	XG10678 	(g24474,g23620);
	not 	XG10679 	(g24463,g23578);
	and 	XG10680 	(g26020,g25034,g9559);
	not 	XG10681 	(g26605,g25293);
	and 	XG10682 	(g24551,g23331,g17148);
	or 	XG10683 	(g25940,g22218,g24415);
	and 	XG10684 	(g25802,g24586,g8106);
	and 	XG10685 	(g26023,g25036,g9528);
	and 	XG10686 	(g25966,g24985,g9364);
	not 	XG10687 	(g26518,g25233);
	and 	XG10688 	(g25969,g24987,g9310);
	nand 	XG10689 	(g20161,g14625,g17670,g17706,g17732);
	and 	XG10690 	(g25876,g24667,g3470);
	and 	XG10691 	(g25879,g24683,g11135);
	and 	XG10692 	(g25875,g24809,g8390);
	or 	XG10693 	(g25943,g22299,g24423);
	and 	XG10694 	(g26323,g25273,g10262);
	not 	XG10695 	(g26548,g25255);
	nor 	XG10696 	(g25932,g24528,g7680);
	and 	XG10697 	(g26815,g24528,g4108);
	or 	XG10698 	(g26089,g22534,g24501);
	not 	XG10699 	(I24128,g23009);
	and 	XG10700 	(g26823,g13106,g24401);
	not 	XG10701 	(g26830,g24411);
	not 	XG10702 	(g25892,g24528);
	nand 	XG10703 	(g20371,g16660,g16694,g14088,g16956);
	nand 	XG10704 	(g21350,g13108,g15735,g15742,g15751);
	or 	XG10705 	(g25935,g22208,g24402);
	nand 	XG10706 	(g21509,g17608,g17647,g14898,g17820);
	not 	XG10707 	(I25028,g24484);
	or 	XG10708 	(g25945,g22307,g24427);
	and 	XG10709 	(g23551,g18948,g10793);
	or 	XG10710 	(g23997,g17191,g20602);
	and 	XG10711 	(g25804,g24587,g8069);
	and 	XG10712 	(g25852,g24411,g4593);
	and 	XG10713 	(g25818,g24605,g8124);
	nand 	XG10714 	(g26752,g25189,g9397);
	and 	XG10715 	(g23475,g8971,g19070);
	and 	XG10716 	(g25788,g24579,g8010);
	and 	XG10717 	(g24774,g23614,g718);
	nand 	XG10718 	(g21603,g17689,g17723,g14987,g17872);
	and 	XG10719 	(g25990,g25017,g9461);
	nand 	XG10720 	(g26208,g24751,g7975);
	nand 	XG10721 	(I23118,g417,g20076);
	and 	XG10722 	(g24719,g23530,g681);
	and 	XG10723 	(g26096,g25268,g9733);
	and 	XG10724 	(g25833,g24626,g8228);
	and 	XG10725 	(g25880,g24814,g8443);
	and 	XG10726 	(g26780,g24437,g4098);
	not 	XG10727 	(g26869,g24842);
	and 	XG10728 	(g26145,g25131,g11962);
	and 	XG10729 	(g26121,g25111,g6167);
	nor 	XG10730 	(g24453,g22325,g7446);
	and 	XG10731 	(g25063,g22325,g13078);
	and 	XG10732 	(g24630,g14149,g23255);
	nand 	XG10733 	(g26666,g25144,g9229);
	and 	XG10734 	(g25801,g24585,g8097);
	not 	XG10735 	(g26054,g24804);
	nor 	XG10736 	(g25521,g14645,g23955);
	and 	XG10737 	(g24786,g23654,g661);
	and 	XG10738 	(g24762,g23573,g655);
	nor 	XG10739 	(g25501,g14645,g23918);
	nor 	XG10740 	(g25247,g14645,g23763);
	nor 	XG10741 	(g26162,g24751,g23052);
	and 	XG10742 	(g25565,g22660,g13013);
	and 	XG10743 	(g26146,g25334,g9892);
	and 	XG10744 	(g25987,g25015,g9501);
	not 	XG10745 	(g26575,g25268);
	nor 	XG10746 	(g25446,g14645,g23686);
	nor 	XG10747 	(g25447,g14645,g23883);
	nor 	XG10748 	(g24391,g14645,g22190);
	and 	XG10749 	(g24676,g23782,g2748);
	nor 	XG10750 	(g25317,g23782,g9766);
	and 	XG10751 	(g24700,g23512,g645);
	and 	XG10752 	(g25832,g24625,g8219);
	not 	XG10753 	(g26093,g24814);
	and 	XG10754 	(g24651,g23472,g2741);
	and 	XG10755 	(g24745,g23550,g650);
	and 	XG10756 	(g24674,g23496,g446);
	nor 	XG10757 	(g26686,g25189,g23678);
	nor 	XG10758 	(g26625,g25144,g23560);
	and 	XG10759 	(g25871,g24804,g8334);
	nand 	XG10760 	(g26255,g24779,g8075);
	nor 	XG10761 	(g26209,g24779,g23124);
	nand 	XG10762 	(g26714,g25175,g9316);
	nor 	XG10763 	(g26667,g25175,g23642);
	and 	XG10764 	(g21997,g19074,g5619);
	and 	XG10765 	(g21770,g20785,g3251);
	not 	XG10766 	(g22881,I22096);
	and 	XG10767 	(g21798,g20924,g3522);
	and 	XG10768 	(g21948,g18997,g5260);
	and 	XG10769 	(g21782,g20391,g3416);
	not 	XG10770 	(g21905,I21486);
	and 	XG10771 	(g21763,g20785,g3223);
	and 	XG10772 	(g21967,g21514,g5456);
	and 	XG10773 	(g21721,g21037,g385);
	and 	XG10774 	(g25374,I24527,g23789,g5366);
	and 	XG10775 	(g21952,g21514,g5366);
	and 	XG10776 	(g21780,g20391,g3391);
	and 	XG10777 	(g21758,g20785,g3191);
	and 	XG10778 	(g21839,g20453,g3763);
	and 	XG10779 	(g21757,g20785,g3187);
	and 	XG10780 	(g21747,g20330,g3061);
	and 	XG10781 	(g21971,g21514,g5417);
	and 	XG10782 	(g22085,g19210,g6295);
	and 	XG10783 	(g21951,g18997,g5272);
	and 	XG10784 	(g21883,g19801,g4141);
	and 	XG10785 	(g21819,g20924,g3614);
	and 	XG10786 	(g21991,g19074,g5595);
	and 	XG10787 	(g21756,g20785,g3211);
	and 	XG10788 	(g21850,g21070,g3893);
	and 	XG10789 	(g22135,g19277,g6657);
	and 	XG10790 	(g21910,g21468,g5016);
	and 	XG10791 	(g21704,g20283,g164);
	and 	XG10792 	(g21838,g20453,g3747);
	and 	XG10793 	(g22017,g21562,g5763);
	and 	XG10794 	(g21911,g21468,g5046);
	and 	XG10795 	(g21936,g18997,g5200);
	and 	XG10796 	(g21882,g19801,g4057);
	and 	XG10797 	(g22049,g21611,g6082);
	and 	XG10798 	(g21737,g20330,g3068);
	and 	XG10799 	(g21862,g21070,g3953);
	not 	XG10800 	(g21722,I21285);
	and 	XG10801 	(g21822,g20453,g3727);
	and 	XG10802 	(g22086,g19210,g6299);
	and 	XG10803 	(g21928,g18997,g5170);
	not 	XG10804 	(g22904,I22111);
	and 	XG10805 	(I24674,g24021,g24020,g24019,g19919);
	and 	XG10806 	(g24897,I24064,g23223,g3401);
	and 	XG10807 	(g21788,g20391,g3401);
	and 	XG10808 	(g21992,g19074,g5599);
	and 	XG10809 	(g22125,g19277,g6617);
	not 	XG10810 	(g21725,I21294);
	and 	XG10811 	(g22028,g19147,g5893);
	and 	XG10812 	(g22054,g21611,g6120);
	and 	XG10813 	(I24695,g24053,g24052,g24051,g24050);
	and 	XG10814 	(I24700,g24060,g24059,g24058,g24057);
	and 	XG10815 	(I24705,g24067,g24066,g24065,g24064);
	not 	XG10816 	(g23444,I22561);
	and 	XG10817 	(I24710,g24074,g24073,g24072,g24071);
	and 	XG10818 	(I24689,g24042,g24041,g24040,g20841);
	and 	XG10819 	(g21965,g21514,g15149);
	and 	XG10820 	(g21771,g20785,g3255);
	and 	XG10821 	(g25488,I24603,g23865,g6404);
	and 	XG10822 	(g22090,g18833,g6404);
	and 	XG10823 	(g22113,g19277,g6561);
	and 	XG10824 	(g22016,g21562,g5747);
	and 	XG10825 	(g21848,g21070,g3913);
	and 	XG10826 	(g21754,g20785,g3195);
	not 	XG10827 	(g22980,I22153);
	and 	XG10828 	(I24684,g24035,g24034,g24033,g20014);
	and 	XG10829 	(g21805,g20924,g3550);
	and 	XG10830 	(g22108,g18833,g6439);
	and 	XG10831 	(g22040,g19147,g5953);
	and 	XG10832 	(g21736,g20330,g3065);
	and 	XG10833 	(g22000,g21562,g5727);
	and 	XG10834 	(g21814,g20924,g3594);
	and 	XG10835 	(g21781,g20391,g3408);
	and 	XG10836 	(g21970,g21514,g5401);
	not 	XG10837 	(g22189,I21769);
	and 	XG10838 	(g25578,g24146,g19402);
	and 	XG10839 	(g21720,g21037,g376);
	and 	XG10840 	(g21873,g19801,g6946);
	and 	XG10841 	(g21922,g21468,g5112);
	and 	XG10842 	(g21761,g20785,g3215);
	and 	XG10843 	(g21918,g21468,g5097);
	and 	XG10844 	(g21945,g18997,g5248);
	and 	XG10845 	(g21772,g20785,g3259);
	and 	XG10846 	(g21760,g20785,g3207);
	and 	XG10847 	(g21890,g19801,g4125);
	not 	XG10848 	(g23481,I22604);
	and 	XG10849 	(I27504,g24080,g24079,g24078,g24077);
	and 	XG10850 	(I27509,g24087,g24086,g24085,g24084);
	and 	XG10851 	(I27514,g24094,g24093,g24092,g24091);
	and 	XG10852 	(I26531,g24102,g24101,g24100,g24099);
	and 	XG10853 	(I27533,g24127,g24126,g24125,g21143);
	and 	XG10854 	(g22026,g19147,g5913);
	not 	XG10855 	(g23480,I22601);
	and 	XG10856 	(I24675,g24025,g24024,g24023,g24022);
	and 	XG10857 	(I24680,g24032,g24031,g24030,g24029);
	and 	XG10858 	(I24685,g24039,g24038,g24037,g24036);
	and 	XG10859 	(I24690,g24046,g24045,g24044,g24043);
	and 	XG10860 	(I24699,g24056,g24055,g24054,g21127);
	and 	XG10861 	(g21759,g20785,g3199);
	and 	XG10862 	(g21907,g21468,g5033);
	and 	XG10863 	(g21876,g19801,g4119);
	and 	XG10864 	(g21940,g18997,g5228);
	and 	XG10865 	(g22102,g18833,g6479);
	or 	XG10866 	(g24577,g22531,g2856);
	or 	XG10867 	(g24705,g23267,g2890);
	and 	XG10868 	(g21818,g20924,g3610);
	and 	XG10869 	(g22117,g19277,g6597);
	and 	XG10870 	(g22119,g19277,g6581);
	and 	XG10871 	(g21776,g20391,g3376);
	and 	XG10872 	(g22122,g19277,g6601);
	and 	XG10873 	(g21785,g20391,g3431);
	and 	XG10874 	(g21762,g20785,g3219);
	and 	XG10875 	(g21718,g21037,g370);
	and 	XG10876 	(g21859,g21070,g3941);
	not 	XG10877 	(g22207,I21787);
	and 	XG10878 	(g21740,g20330,g3085);
	and 	XG10879 	(g21878,g19801,g4129);
	and 	XG10880 	(g22114,g19277,g6565);
	and 	XG10881 	(g22096,g18833,g6434);
	and 	XG10882 	(g22053,g21611,g6116);
	and 	XG10883 	(g21874,g19801,g4112);
	and 	XG10884 	(g21953,g21514,g5377);
	not 	XG10885 	(g22159,I21744);
	and 	XG10886 	(g25581,g24150,g19338);
	and 	XG10887 	(g21854,g21070,g3921);
	and 	XG10888 	(g21913,g21468,g5069);
	and 	XG10889 	(g22087,g19210,g6303);
	not 	XG10890 	(g23430,I22547);
	and 	XG10891 	(I27518,g24106,g24105,g24104,g20720);
	and 	XG10892 	(g22129,g19277,g6633);
	and 	XG10893 	(g21925,g21468,g5073);
	and 	XG10894 	(g22097,g18833,g6451);
	and 	XG10895 	(g22093,g18833,g6423);
	or 	XG10896 	(g24264,g18559,g22310);
	and 	XG10897 	(g21717,g21037,g15051);
	and 	XG10898 	(g21929,g18997,g5176);
	and 	XG10899 	(g21946,g18997,g5252);
	and 	XG10900 	(g22037,g19147,g5941);
	and 	XG10901 	(g21885,g19801,g4122);
	not 	XG10902 	(g23457,I22580);
	and 	XG10903 	(I24694,g24049,g24048,g24047,g20982);
	and 	XG10904 	(g21926,g18997,g15147);
	and 	XG10905 	(g21823,g20453,g3731);
	and 	XG10906 	(g21748,g20785,g15089);
	or 	XG10907 	(g24363,g22138,g7831);
	and 	XG10908 	(g22115,g19277,g6573);
	and 	XG10909 	(g21920,g21468,g5062);
	and 	XG10910 	(g25411,I24546,g23764,g5062);
	and 	XG10911 	(g22101,g18833,g6474);
	and 	XG10912 	(g21703,g20283,g146);
	and 	XG10913 	(g22032,g19147,g5921);
	and 	XG10914 	(g22107,g18833,g6411);
	and 	XG10915 	(g21813,g20924,g3590);
	and 	XG10916 	(g25459,I24582,g23844,g6058);
	and 	XG10917 	(g22044,g21611,g6058);
	and 	XG10918 	(g21933,g18997,g5212);
	and 	XG10919 	(g22120,g19277,g6585);
	and 	XG10920 	(g22118,g19277,g6605);
	not 	XG10921 	(g23445,I22564);
	and 	XG10922 	(I27523,g24113,g24112,g24111,g20857);
	and 	XG10923 	(g22001,g21562,g5731);
	and 	XG10924 	(g21860,g21070,g3945);
	and 	XG10925 	(g22077,g19210,g6263);
	or 	XG10926 	(g24965,g23825,g22667);
	and 	XG10927 	(g21984,g19074,g5563);
	and 	XG10928 	(g22062,g21611,g6093);
	not 	XG10929 	(g23495,I22622);
	and 	XG10930 	(I27538,g24134,g24133,g24132,g21209);
	and 	XG10931 	(g21855,g21070,g3925);
	and 	XG10932 	(g21942,g18997,g5236);
	and 	XG10933 	(g21800,g20924,g3546);
	and 	XG10934 	(g22056,g21611,g6133);
	and 	XG10935 	(g21732,g20330,g3004);
	and 	XG10936 	(g22109,g18833,g6455);
	and 	XG10937 	(g22100,g18833,g6466);
	and 	XG10938 	(g22116,g19277,g6589);
	and 	XG10939 	(g21974,g19074,g5517);
	and 	XG10940 	(g22123,g19277,g6609);
	and 	XG10941 	(g21705,g20283,g209);
	and 	XG10942 	(g21944,g18997,g5244);
	and 	XG10943 	(g22038,g19147,g5945);
	and 	XG10944 	(g21861,g21070,g3949);
	and 	XG10945 	(g22075,g19210,g6247);
	and 	XG10946 	(g22095,g18833,g6428);
	and 	XG10947 	(g21831,g20453,g3782);
	and 	XG10948 	(g21982,g19074,g5547);
	not 	XG10949 	(g21724,I21291);
	and 	XG10950 	(g22065,g19210,g6203);
	and 	XG10951 	(g21939,g18997,g5224);
	and 	XG10952 	(g22033,g19147,g5925);
	and 	XG10953 	(g21856,g21070,g3929);
	and 	XG10954 	(g22069,g19210,g6227);
	and 	XG10955 	(g22091,g18833,g6415);
	and 	XG10956 	(g21976,g19074,g5527);
	and 	XG10957 	(g22098,g18833,g6459);
	and 	XG10958 	(g22082,g19210,g6283);
	and 	XG10959 	(g21988,g19074,g5583);
	and 	XG10960 	(g21881,g19801,g4064);
	and 	XG10961 	(g21993,g19074,g5603);
	and 	XG10962 	(g21916,g21468,g5084);
	and 	XG10963 	(g22051,g21611,g6105);
	and 	XG10964 	(g22103,g18833,g15164);
	and 	XG10965 	(g22039,g19147,g5949);
	and 	XG10966 	(g22009,g21562,g5782);
	and 	XG10967 	(g21858,g21070,g3937);
	and 	XG10968 	(g21867,g19801,g4082);
	and 	XG10969 	(g22034,g19147,g5929);
	and 	XG10970 	(g22048,g21611,g6052);
	and 	XG10971 	(g22092,g18833,g6419);
	and 	XG10972 	(g21707,g20283,g191);
	and 	XG10973 	(g22058,g21611,g6098);
	and 	XG10974 	(g25507,I24616,g23844,g6098);
	and 	XG10975 	(g21733,g20330,g3034);
	and 	XG10976 	(g21738,g20330,g3072);
	and 	XG10977 	(g21957,g21514,g5390);
	and 	XG10978 	(g22063,g21611,g6109);
	and 	XG10979 	(g21744,g20330,g3103);
	and 	XG10980 	(g22036,g19147,g5937);
	and 	XG10981 	(g21789,g20391,g3451);
	and 	XG10982 	(g21774,g20391,g3361);
	and 	XG10983 	(g24858,I24030,g23223,g3361);
	and 	XG10984 	(g21750,g20785,g3161);
	and 	XG10985 	(g21709,g20283,g283);
	and 	XG10986 	(g21784,g20391,g3423);
	not 	XG10987 	(g21723,I21288);
	and 	XG10988 	(g21719,g21037,g358);
	and 	XG10989 	(g21959,g21514,g5413);
	and 	XG10990 	(g21841,g21070,g3857);
	and 	XG10991 	(g22134,g19277,g6653);
	not 	XG10992 	(g22927,I22128);
	nor 	XG10993 	(g24018,I23163,I23162);
	and 	XG10994 	(g21842,g21070,g3863);
	and 	XG10995 	(g21739,g20330,g3080);
	and 	XG10996 	(g21943,g18997,g5240);
	and 	XG10997 	(g25479,g9917,g22646);
	and 	XG10998 	(g21791,g20391,g3368);
	and 	XG10999 	(g21934,g18997,g5220);
	and 	XG11000 	(g21710,g20283,g287);
	not 	XG11001 	(g22928,I22131);
	and 	XG11002 	(g21821,g20453,g3723);
	and 	XG11003 	(g21802,g20924,g3562);
	and 	XG11004 	(g22019,g19147,g5857);
	and 	XG11005 	(g25518,I24625,g23865,g6444);
	and 	XG11006 	(g22104,g18833,g6444);
	and 	XG11007 	(g22124,g19277,g6613);
	and 	XG11008 	(g21773,g20785,g3263);
	and 	XG11009 	(g21729,g20330,g3021);
	and 	XG11010 	(g22020,g19147,g5863);
	and 	XG11011 	(g21915,g21468,g5080);
	not 	XG11012 	(g23511,I22640);
	and 	XG11013 	(g21708,g20283,g15049);
	and 	XG11014 	(g22047,g21611,g6077);
	or 	XG11015 	(g24212,g18155,g23280);
	and 	XG11016 	(g21716,g20283,g301);
	and 	XG11017 	(g21803,g20924,g3538);
	and 	XG11018 	(g21792,g20391,g3396);
	and 	XG11019 	(g21830,g20453,g3774);
	and 	XG11020 	(g21713,g20283,g298);
	and 	XG11021 	(g21964,g21514,g5441);
	and 	XG11022 	(g21909,g21468,g5041);
	and 	XG11023 	(g21875,g19801,g4116);
	not 	XG11024 	(g22905,I22114);
	and 	XG11025 	(g21866,g19801,g4072);
	not 	XG11026 	(g23458,I22583);
	and 	XG11027 	(g21999,g21562,g5723);
	and 	XG11028 	(g25408,g9772,g22682);
	and 	XG11029 	(g21769,g20785,g3247);
	and 	XG11030 	(g21960,g21514,g5421);
	and 	XG11031 	(g21954,g21514,g5381);
	and 	XG11032 	(g21947,g18997,g5256);
	and 	XG11033 	(g22066,g19210,g6209);
	and 	XG11034 	(g21755,g20785,g3203);
	and 	XG11035 	(g21764,g20785,g3227);
	and 	XG11036 	(g21958,g21514,g5396);
	and 	XG11037 	(g21935,g18997,g5196);
	and 	XG11038 	(g22008,g21562,g5774);
	and 	XG11039 	(g22079,g19210,g6271);
	and 	XG11040 	(g21811,g20924,g3582);
	and 	XG11041 	(g21828,g20453,g3767);
	and 	XG11042 	(g21810,g20924,g3578);
	and 	XG11043 	(g21985,g19074,g5571);
	and 	XG11044 	(g21816,g20924,g3602);
	and 	XG11045 	(g21746,g20330,g3045);
	and 	XG11046 	(g22131,g19277,g6641);
	and 	XG11047 	(g22121,g19277,g6593);
	and 	XG11048 	(g21962,g21514,g5428);
	and 	XG11049 	(g22105,g18833,g6494);
	and 	XG11050 	(g21938,g18997,g5216);
	and 	XG11051 	(g21931,g18997,g5188);
	and 	XG11052 	(g22052,g21611,g6113);
	and 	XG11053 	(g21730,g20330,g3025);
	and 	XG11054 	(g21846,g21070,g3897);
	and 	XG11055 	(g22126,g19277,g6621);
	and 	XG11056 	(g21845,g21070,g3881);
	and 	XG11057 	(g21779,g20391,g3385);
	and 	XG11058 	(g22112,g19277,g6555);
	and 	XG11059 	(g21700,g20283,g150);
	and 	XG11060 	(g22073,g19210,g6235);
	and 	XG11061 	(g21783,g20391,g3419);
	and 	XG11062 	(g21977,g19074,g5535);
	and 	XG11063 	(g22006,g21562,g5767);
	and 	XG11064 	(g21968,g21514,g5459);
	and 	XG11065 	(g21969,g21514,g5373);
	and 	XG11066 	(g21972,g19074,g15152);
	and 	XG11067 	(g21715,g20283,g160);
	and 	XG11068 	(g22060,g21611,g6151);
	and 	XG11069 	(g21870,g19801,g4093);
	and 	XG11070 	(g21863,g21070,g3957);
	and 	XG11071 	(g21827,g20453,g3759);
	and 	XG11072 	(g21840,g21070,g15099);
	and 	XG11073 	(g21966,g21514,g5406);
	and 	XG11074 	(g25453,I24576,g23789,g5406);
	and 	XG11075 	(g21787,g20391,g15091);
	and 	XG11076 	(g21888,g19801,g4165);
	and 	XG11077 	(g22024,g19147,g5897);
	and 	XG11078 	(g21832,g20453,g3787);
	and 	XG11079 	(g21752,g20785,g3171);
	and 	XG11080 	(g21731,g20330,g3029);
	and 	XG11081 	(g22023,g19147,g5881);
	and 	XG11082 	(g21955,g21514,g5385);
	and 	XG11083 	(g21833,g20453,g15096);
	and 	XG11084 	(g21824,g20453,g3706);
	and 	XG11085 	(g21793,g20391,g3412);
	and 	XG11086 	(g21871,g19801,g4108);
	and 	XG11087 	(g21912,g21468,g5052);
	not 	XG11088 	(g21903,I21480);
	and 	XG11089 	(g21950,g18997,g5268);
	and 	XG11090 	(g21829,g20453,g3770);
	and 	XG11091 	(g22074,g19210,g6239);
	and 	XG11092 	(g21790,g20391,g3454);
	and 	XG11093 	(g22089,g19210,g6311);
	and 	XG11094 	(g22080,g19210,g6275);
	and 	XG11095 	(g21853,g21070,g3917);
	and 	XG11096 	(g24908,I24075,g23239,g3752);
	and 	XG11097 	(g21834,g20453,g3752);
	and 	XG11098 	(g21986,g19074,g5575);
	and 	XG11099 	(g21837,g20453,g3719);
	and 	XG11100 	(g21843,g21070,g3869);
	and 	XG11101 	(g22041,g19147,g5957);
	and 	XG11102 	(g21844,g21070,g3873);
	and 	XG11103 	(g22005,g21562,g5759);
	and 	XG11104 	(g22132,g19277,g6645);
	and 	XG11105 	(g22018,g19147,g15157);
	and 	XG11106 	(g21921,g21468,g5109);
	and 	XG11107 	(g21836,g20453,g3805);
	and 	XG11108 	(g21919,g21468,g15144);
	and 	XG11109 	(g21741,g20330,g15086);
	and 	XG11110 	(g22010,g21562,g5787);
	and 	XG11111 	(g21786,g20391,g3436);
	and 	XG11112 	(g21889,g19801,g4169);
	and 	XG11113 	(g21923,g21468,g5029);
	and 	XG11114 	(g22011,g21562,g15154);
	and 	XG11115 	(g22002,g21562,g5706);
	and 	XG11116 	(g22127,g19277,g6625);
	not 	XG11117 	(g22151,I21734);
	and 	XG11118 	(g22007,g21562,g5770);
	and 	XG11119 	(g21864,g21070,g3961);
	and 	XG11120 	(g21869,g19801,g4087);
	and 	XG11121 	(g22111,g19277,g6549);
	and 	XG11122 	(g21701,g20283,g153);
	and 	XG11123 	(g21927,g18997,g5164);
	and 	XG11124 	(g24887,I24054,g23239,g3712);
	and 	XG11125 	(g21820,g20453,g3712);
	not 	XG11126 	(g21726,I21297);
	and 	XG11127 	(g22031,g19147,g5917);
	and 	XG11128 	(g22081,g19210,g6279);
	and 	XG11129 	(g25482,I24597,g23816,g5752);
	and 	XG11130 	(g22012,g21562,g5752);
	and 	XG11131 	(g22015,g21562,g5719);
	and 	XG11132 	(g22021,g19147,g5869);
	and 	XG11133 	(g21987,g19074,g5579);
	and 	XG11134 	(g21937,g18997,g5208);
	and 	XG11135 	(g21908,g21468,g5037);
	and 	XG11136 	(g22022,g19147,g5873);
	and 	XG11137 	(g21826,g20453,g3742);
	and 	XG11138 	(g22133,g19277,g6649);
	and 	XG11139 	(g22059,g21611,g6148);
	and 	XG11140 	(g21765,g20785,g3231);
	and 	XG11141 	(g21906,g21468,g5022);
	and 	XG11142 	(g25328,I24505,g23764,g5022);
	and 	XG11143 	(g22014,g21562,g5805);
	or 	XG11144 	(g24653,g22585,g2848);
	and 	XG11145 	(g21699,g20283,g142);
	and 	XG11146 	(g21963,g21514,g5436);
	and 	XG11147 	(g21872,g19801,g4098);
	or 	XG11148 	(g25010,g2932,g23267);
	and 	XG11149 	(g22128,g19277,g6629);
	and 	XG11150 	(g22055,g21611,g6128);
	and 	XG11151 	(g21849,g21070,g3889);
	and 	XG11152 	(g22070,g19210,g6243);
	and 	XG11153 	(g22042,g19147,g5961);
	and 	XG11154 	(g21825,g20453,g3736);
	and 	XG11155 	(g21981,g19074,g5543);
	and 	XG11156 	(g25417,I24552,g23816,g5712);
	and 	XG11157 	(g21998,g21562,g5712);
	and 	XG11158 	(g21809,g20924,g3574);
	and 	XG11159 	(g21702,g20283,g157);
	and 	XG11160 	(g22071,g19210,g6251);
	and 	XG11161 	(g21851,g21070,g3901);
	and 	XG11162 	(g21806,g20924,g3558);
	and 	XG11163 	(g22004,g21562,g5742);
	and 	XG11164 	(g21978,g19074,g5551);
	and 	XG11165 	(g21835,g20453,g3802);
	and 	XG11166 	(g22088,g19210,g6307);
	and 	XG11167 	(g22130,g19277,g6637);
	and 	XG11168 	(g21975,g19074,g5523);
	and 	XG11169 	(g21914,g21468,g5077);
	not 	XG11170 	(g23494,I22619);
	and 	XG11171 	(g21961,g21514,g5424);
	and 	XG11172 	(g21877,g19801,g6888);
	and 	XG11173 	(g21753,g20785,g3179);
	and 	XG11174 	(g22027,g19147,g5889);
	and 	XG11175 	(g22110,g19277,g15167);
	and 	XG11176 	(g22003,g21562,g5736);
	and 	XG11177 	(g24881,I24048,g23211,g3050);
	and 	XG11178 	(g21742,g20330,g3050);
	and 	XG11179 	(g21706,g20283,g222);
	and 	XG11180 	(g21857,g21070,g3933);
	and 	XG11181 	(g21865,g21070,g3965);
	and 	XG11182 	(g21917,g21468,g5092);
	and 	XG11183 	(g21880,g19801,g4135);
	and 	XG11184 	(g21797,g20924,g3518);
	and 	XG11185 	(g21973,g19074,g5511);
	and 	XG11186 	(g22029,g19147,g5901);
	and 	XG11187 	(g22013,g21562,g5802);
	not 	XG11188 	(g21904,I21483);
	and 	XG11189 	(g22094,g18833,g6398);
	and 	XG11190 	(g21807,g20924,g3566);
	and 	XG11191 	(g21766,g20785,g3235);
	and 	XG11192 	(g21995,g19074,g5611);
	and 	XG11193 	(g21775,g20391,g3372);
	and 	XG11194 	(g21728,g20330,g3010);
	and 	XG11195 	(g24843,I24015,g23211,g3010);
	and 	XG11196 	(g21884,g19801,g4104);
	and 	XG11197 	(g21799,g20924,g3530);
	or 	XG11198 	(g24213,g18186,g23220);
	and 	XG11199 	(g22035,g19147,g5933);
	and 	XG11200 	(g21956,g21514,g5360);
	and 	XG11201 	(g21949,g18997,g5264);
	and 	XG11202 	(g22043,g19147,g5965);
	and 	XG11203 	(g21794,g20924,g15094);
	and 	XG11204 	(g22078,g19210,g6267);
	not 	XG11205 	(g21902,I21477);
	and 	XG11206 	(g21734,g20330,g3040);
	and 	XG11207 	(g21980,g19074,g5567);
	and 	XG11208 	(g22106,g18833,g6497);
	and 	XG11209 	(g21743,g20330,g3100);
	and 	XG11210 	(g22076,g19210,g6255);
	and 	XG11211 	(g21847,g21070,g3905);
	and 	XG11212 	(g21868,g19801,g4076);
	and 	XG11213 	(g21983,g19074,g5555);
	and 	XG11214 	(g21887,g19801,g15101);
	and 	XG11215 	(g21777,g20391,g3380);
	and 	XG11216 	(g22064,g19210,g15162);
	and 	XG11217 	(g21767,g20785,g3239);
	and 	XG11218 	(g21714,g20283,g278);
	and 	XG11219 	(g22061,g21611,g6065);
	and 	XG11220 	(g21795,g20924,g3506);
	and 	XG11221 	(g22057,g21611,g15159);
	and 	XG11222 	(g21886,g19801,g4153);
	and 	XG11223 	(g21879,g19801,g4132);
	and 	XG11224 	(g21808,g20924,g3570);
	and 	XG11225 	(g21711,g20283,g291);
	and 	XG11226 	(g21812,g20924,g3586);
	and 	XG11227 	(g22067,g19210,g6215);
	and 	XG11228 	(g21817,g20924,g3606);
	and 	XG11229 	(g21932,g18997,g5204);
	and 	XG11230 	(g22050,g21611,g6088);
	and 	XG11231 	(g22025,g19147,g5905);
	and 	XG11232 	(g22072,g19210,g6259);
	and 	XG11233 	(g21852,g21070,g3909);
	and 	XG11234 	(g21979,g19074,g5559);
	and 	XG11235 	(g21712,g20283,g294);
	and 	XG11236 	(g22084,g19210,g6291);
	and 	XG11237 	(g21815,g20924,g3598);
	and 	XG11238 	(g21990,g19074,g5591);
	and 	XG11239 	(g21930,g18997,g5180);
	and 	XG11240 	(g22083,g19210,g6287);
	and 	XG11241 	(g21735,g20330,g3057);
	and 	XG11242 	(g21996,g19074,g5615);
	and 	XG11243 	(g21751,g20785,g3167);
	and 	XG11244 	(g21989,g19074,g5587);
	and 	XG11245 	(g22045,g21611,g6069);
	and 	XG11246 	(g21994,g19074,g5607);
	and 	XG11247 	(g22046,g21611,g6073);
	and 	XG11248 	(g21778,g20391,g3355);
	and 	XG11249 	(g21749,g20785,g3155);
	and 	XG11250 	(g21796,g20924,g3512);
	and 	XG11251 	(g22068,g19210,g6219);
	and 	XG11252 	(g21801,g20924,g3554);
	and 	XG11253 	(g22030,g19147,g5909);
	and 	XG11254 	(g21941,g18997,g5232);
	and 	XG11255 	(g21804,g20924,g3542);
	and 	XG11256 	(g21768,g20785,g3243);
	and 	XG11257 	(g21745,g20330,g3017);
	and 	XG11258 	(g22099,g18833,g6462);
	and 	XG11259 	(g21924,g21468,g5057);
	not 	XG11260 	(g22202,I21784);
	not 	XG11261 	(g22409,I21860);
	not 	XG11262 	(g23320,I22419);
	not 	XG11263 	(g23232,I22331);
	not 	XG11264 	(g23395,I22502);
	not 	XG11265 	(g23263,I22366);
	not 	XG11266 	(g23427,I22542);
	not 	XG11267 	(g23361,I22464);
	not 	XG11268 	(g23299,I22400);
	not 	XG11269 	(g22360,I21849);
	not 	XG11270 	(g22182,I21766);
	not 	XG11271 	(g23414,I22525);
	not 	XG11272 	(g23347,I22444);
	not 	XG11273 	(g23362,I22467);
	not 	XG11274 	(g23322,I22425);
	not 	XG11275 	(g22658,I21969);
	nand 	XG11276 	(g24362,g22136,g21370);
	not 	XG11277 	(g23385,I22488);
	not 	XG11278 	(g22721,I22028);
	not 	XG11279 	(g23450,I22571);
	not 	XG11280 	(g23277,I22380);
	not 	XG11281 	(g22683,I22000);
	not 	XG11282 	(g23359,I22458);
	not 	XG11283 	(g23403,I22512);
	not 	XG11284 	(g22647,I21959);
	not 	XG11285 	(g23360,I22461);
	not 	XG11286 	(g23394,I22499);
	not 	XG11287 	(g23321,I22422);
	not 	XG11288 	(g22763,I22046);
	not 	XG11289 	(g23426,I22539);
	not 	XG11290 	(g23555,I22692);
	not 	XG11291 	(g22194,I21776);
	not 	XG11292 	(g22300,I21815);
	not 	XG11293 	(g22173,I21757);
	not 	XG11294 	(g22220,I21802);
	not 	XG11295 	(g22210,I21792);
	not 	XG11296 	(g23534,I22665);
	not 	XG11297 	(g23384,I22485);
	not 	XG11298 	(g23582,I22729);
	not 	XG11299 	(g23378,g21070);
	not 	XG11300 	(g23228,g21070);
	not 	XG11301 	(g23356,g21070);
	not 	XG11302 	(g23249,g21070);
	not 	XG11303 	(g23274,g21070);
	not 	XG11304 	(g23517,g21070);
	not 	XG11305 	(g23340,g21070);
	not 	XG11306 	(g23242,g21070);
	not 	XG11307 	(g23502,g21070);
	not 	XG11308 	(g23243,g21070);
	not 	XG11309 	(g23339,g21070);
	not 	XG11310 	(g23250,g21070);
	not 	XG11311 	(g23376,g21070);
	not 	XG11312 	(g23377,g21070);
	not 	XG11313 	(g23355,g21070);
	not 	XG11314 	(g23388,g21070);
	not 	XG11315 	(g23291,g21070);
	not 	XG11316 	(g23273,g21070);
	not 	XG11317 	(g23539,g21070);
	not 	XG11318 	(g23312,g21070);
	not 	XG11319 	(g23585,g21070);
	not 	XG11320 	(g23518,g21070);
	not 	XG11321 	(g23313,g21070);
	not 	XG11322 	(g23559,g21070);
	not 	XG11323 	(g23260,g21070);
	not 	XG11324 	(g23259,g21070);
	not 	XG11325 	(g23057,g20453);
	not 	XG11326 	(g23429,g20453);
	not 	XG11327 	(g22868,g20453);
	not 	XG11328 	(g22989,g20453);
	not 	XG11329 	(g22856,g20453);
	not 	XG11330 	(g22999,g20453);
	not 	XG11331 	(g23000,g20453);
	not 	XG11332 	(g23338,g20453);
	not 	XG11333 	(g22884,g20453);
	not 	XG11334 	(g23354,g20453);
	not 	XG11335 	(g23058,g20453);
	not 	XG11336 	(g23059,g20453);
	not 	XG11337 	(g22979,g20453);
	not 	XG11338 	(g23029,g20453);
	not 	XG11339 	(g23138,g20453);
	not 	XG11340 	(g23030,g20453);
	not 	XG11341 	(g23016,g20453);
	not 	XG11342 	(g22906,g20453);
	not 	XG11343 	(g23017,g20453);
	not 	XG11344 	(g22907,g20453);
	not 	XG11345 	(g23448,g21611);
	not 	XG11346 	(g23945,g21611);
	not 	XG11347 	(g23509,g21611);
	not 	XG11348 	(g23607,g21611);
	not 	XG11349 	(g23422,g21611);
	not 	XG11350 	(g23493,g21611);
	not 	XG11351 	(g24013,g21611);
	not 	XG11352 	(g23568,g21611);
	not 	XG11353 	(g23569,g21611);
	not 	XG11354 	(g23965,g21611);
	not 	XG11355 	(g23526,g21611);
	not 	XG11356 	(g23527,g21611);
	not 	XG11357 	(g23546,g21611);
	not 	XG11358 	(g23547,g21611);
	not 	XG11359 	(g23698,g21611);
	not 	XG11360 	(g23434,g21611);
	not 	XG11361 	(g23608,g21611);
	not 	XG11362 	(g23609,g21611);
	not 	XG11363 	(g23460,g21611);
	not 	XG11364 	(g23459,g21611);
	not 	XG11365 	(g23880,g19210);
	not 	XG11366 	(g23896,g19210);
	not 	XG11367 	(g23897,g19210);
	not 	XG11368 	(g22199,g19210);
	not 	XG11369 	(g23847,g19210);
	not 	XG11370 	(g23821,g19210);
	not 	XG11371 	(g23863,g19210);
	not 	XG11372 	(g23983,g19210);
	not 	XG11373 	(g23992,g19210);
	not 	XG11374 	(g23936,g19210);
	not 	XG11375 	(g22179,g19210);
	not 	XG11376 	(g22223,g19210);
	not 	XG11377 	(g22180,g19210);
	not 	XG11378 	(g23946,g19210);
	not 	XG11379 	(g23947,g19210);
	not 	XG11380 	(g23848,g19210);
	not 	XG11381 	(g23935,g19210);
	not 	XG11382 	(g23914,g19210);
	not 	XG11383 	(g23864,g19210);
	not 	XG11384 	(g23984,g19210);
	not 	XG11385 	(g22214,g19210);
	not 	XG11386 	(g23985,g19210);
	not 	XG11387 	(g23966,g19210);
	not 	XG11388 	(g23967,g19210);
	not 	XG11389 	(g23879,g19210);
	not 	XG11390 	(g22170,g19210);
	not 	XG11391 	(I21934,g21273);
	not 	XG11392 	(g23233,g21037);
	not 	XG11393 	(g23264,g21037);
	not 	XG11394 	(g23253,g21037);
	not 	XG11395 	(g23279,g21037);
	not 	XG11396 	(g23301,g21037);
	not 	XG11397 	(I22031,g21387);
	not 	XG11398 	(g23323,g20283);
	not 	XG11399 	(g23128,g20283);
	not 	XG11400 	(g22830,g20283);
	not 	XG11401 	(g23046,g20283);
	not 	XG11402 	(g23152,g20283);
	not 	XG11403 	(g23021,g20283);
	not 	XG11404 	(g22847,g20283);
	not 	XG11405 	(g23278,g20283);
	not 	XG11406 	(g23300,g20283);
	not 	XG11407 	(g22936,g20283);
	not 	XG11408 	(g23061,g20283);
	not 	XG11409 	(g23004,g20283);
	not 	XG11410 	(g23005,g20283);
	not 	XG11411 	(g22898,g20283);
	not 	XG11412 	(g22981,g20283);
	not 	XG11413 	(g23022,g20283);
	not 	XG11414 	(g22935,g20283);
	not 	XG11415 	(g23086,g20283);
	not 	XG11416 	(g23026,g20391);
	not 	XG11417 	(g23027,g20391);
	not 	XG11418 	(g22988,g20391);
	not 	XG11419 	(g22998,g20391);
	not 	XG11420 	(g23014,g20391);
	not 	XG11421 	(g23417,g20391);
	not 	XG11422 	(g23015,g20391);
	not 	XG11423 	(g23335,g20391);
	not 	XG11424 	(g22841,g20391);
	not 	XG11425 	(g23111,g20391);
	not 	XG11426 	(g22975,g20391);
	not 	XG11427 	(g22867,g20391);
	not 	XG11428 	(g22855,g20391);
	not 	XG11429 	(g22987,g20391);
	not 	XG11430 	(g23028,g20391);
	not 	XG11431 	(g22997,g20391);
	not 	XG11432 	(g22926,g20391);
	not 	XG11433 	(g23305,g20391);
	not 	XG11434 	(g22882,g20391);
	not 	XG11435 	(g22883,g20391);
	not 	XG11436 	(g23248,g20924);
	not 	XG11437 	(g23516,g20924);
	not 	XG11438 	(g23351,g20924);
	not 	XG11439 	(g23237,g20924);
	not 	XG11440 	(g23216,g20924);
	not 	XG11441 	(g23306,g20924);
	not 	XG11442 	(g23487,g20924);
	not 	XG11443 	(g23307,g20924);
	not 	XG11444 	(g23257,g20924);
	not 	XG11445 	(g23226,g20924);
	not 	XG11446 	(g23290,g20924);
	not 	XG11447 	(g23227,g20924);
	not 	XG11448 	(g23272,g20924);
	not 	XG11449 	(g23247,g20924);
	not 	XG11450 	(g23500,g20924);
	not 	XG11451 	(g23538,g20924);
	not 	XG11452 	(g23501,g20924);
	not 	XG11453 	(g23238,g20924);
	not 	XG11454 	(g23352,g20924);
	not 	XG11455 	(g23558,g20924);
	not 	XG11456 	(g23289,g20924);
	not 	XG11457 	(g23336,g20924);
	not 	XG11458 	(g23353,g20924);
	not 	XG11459 	(g23337,g20924);
	not 	XG11460 	(g23375,g20924);
	not 	XG11461 	(g23258,g20924);
	not 	XG11462 	(g22455,g19801);
	not 	XG11463 	(g22495,g19801);
	not 	XG11464 	(g22330,g19801);
	not 	XG11465 	(g22528,g19801);
	not 	XG11466 	(g22317,g19801);
	not 	XG11467 	(g22192,g19801);
	not 	XG11468 	(g22635,g19801);
	not 	XG11469 	(g22593,g19801);
	not 	XG11470 	(g22542,g19801);
	not 	XG11471 	(g23001,g19801);
	not 	XG11472 	(g22493,g19801);
	not 	XG11473 	(g23018,g19801);
	not 	XG11474 	(g22543,g19801);
	not 	XG11475 	(g22341,g19801);
	not 	XG11476 	(g22456,g19801);
	not 	XG11477 	(g22526,g19801);
	not 	XG11478 	(g22338,g19801);
	not 	XG11479 	(g22339,g19801);
	not 	XG11480 	(g22520,g19801);
	not 	XG11481 	(g22227,g19801);
	not 	XG11482 	(g22358,g19801);
	not 	XG11483 	(g22519,g19801);
	not 	XG11484 	(g22305,g19801);
	not 	XG11485 	(g23031,g19801);
	not 	XG11486 	(g22494,g19801);
	not 	XG11487 	(g22144,g18997);
	not 	XG11488 	(g23768,g18997);
	not 	XG11489 	(g23787,g18997);
	not 	XG11490 	(g23904,g18997);
	not 	XG11491 	(g23922,g18997);
	not 	XG11492 	(g22153,g18997);
	not 	XG11493 	(g23838,g18997);
	not 	XG11494 	(g23839,g18997);
	not 	XG11495 	(g23923,g18997);
	not 	XG11496 	(g23888,g18997);
	not 	XG11497 	(g23858,g18997);
	not 	XG11498 	(g23767,g18997);
	not 	XG11499 	(g23903,g18997);
	not 	XG11500 	(g23788,g18997);
	not 	XG11501 	(g23812,g18997);
	not 	XG11502 	(g22146,g18997);
	not 	XG11503 	(g22147,g18997);
	not 	XG11504 	(g23813,g18997);
	not 	XG11505 	(g23874,g18997);
	not 	XG11506 	(g23749,g18997);
	not 	XG11507 	(g23875,g18997);
	not 	XG11508 	(g23938,g18997);
	not 	XG11509 	(g22176,g18997);
	not 	XG11510 	(g22166,g18997);
	not 	XG11511 	(g23887,g18997);
	not 	XG11512 	(g23924,g18997);
	not 	XG11513 	(g23504,g21468);
	not 	XG11514 	(g23999,g21468);
	not 	XG11515 	(g23452,g21468);
	not 	XG11516 	(g23390,g21468);
	not 	XG11517 	(g23408,g21468);
	not 	XG11518 	(g23443,g21468);
	not 	XG11519 	(g23503,g21468);
	not 	XG11520 	(g23520,g21468);
	not 	XG11521 	(g23902,g21468);
	not 	XG11522 	(g23521,g21468);
	not 	XG11523 	(g23398,g21468);
	not 	XG11524 	(g23519,g21468);
	not 	XG11525 	(g23476,g21468);
	not 	XG11526 	(g23477,g21468);
	not 	XG11527 	(g23589,g21468);
	not 	XG11528 	(g23418,g21468);
	not 	XG11529 	(g23419,g21468);
	not 	XG11530 	(g23488,g21468);
	not 	XG11531 	(g23489,g21468);
	not 	XG11532 	(g23886,g21468);
	not 	XG11533 	(I21922,g21335);
	not 	XG11534 	(I21810,g20596);
	not 	XG11535 	(g23944,g19147);
	not 	XG11536 	(g22198,g19147);
	not 	XG11537 	(g23929,g19147);
	not 	XG11538 	(g23820,g19147);
	not 	XG11539 	(g23912,g19147);
	not 	XG11540 	(g23862,g19147);
	not 	XG11541 	(g23982,g19147);
	not 	XG11542 	(g23913,g19147);
	not 	XG11543 	(g22213,g19147);
	not 	XG11544 	(g23964,g19147);
	not 	XG11545 	(g23930,g19147);
	not 	XG11546 	(g23877,g19147);
	not 	XG11547 	(g23819,g19147);
	not 	XG11548 	(g23943,g19147);
	not 	XG11549 	(g22178,g19147);
	not 	XG11550 	(g22168,g19147);
	not 	XG11551 	(g22169,g19147);
	not 	XG11552 	(g23895,g19147);
	not 	XG11553 	(g22156,g19147);
	not 	XG11554 	(g23861,g19147);
	not 	XG11555 	(g23794,g19147);
	not 	XG11556 	(g23962,g19147);
	not 	XG11557 	(g23963,g19147);
	not 	XG11558 	(g23842,g19147);
	not 	XG11559 	(g23878,g19147);
	not 	XG11560 	(g23843,g19147);
	not 	XG11561 	(g23433,g21562);
	not 	XG11562 	(g23928,g21562);
	not 	XG11563 	(g23508,g21562);
	not 	XG11564 	(g23492,g21562);
	not 	XG11565 	(g23565,g21562);
	not 	XG11566 	(g23479,g21562);
	not 	XG11567 	(g23410,g21562);
	not 	XG11568 	(g23942,g21562);
	not 	XG11569 	(g24010,g21562);
	not 	XG11570 	(g23446,g21562);
	not 	XG11571 	(g23447,g21562);
	not 	XG11572 	(g23421,g21562);
	not 	XG11573 	(g23507,g21562);
	not 	XG11574 	(g23566,g21562);
	not 	XG11575 	(g23567,g21562);
	not 	XG11576 	(g23665,g21562);
	not 	XG11577 	(g23524,g21562);
	not 	XG11578 	(g23544,g21562);
	not 	XG11579 	(g23525,g21562);
	not 	XG11580 	(g23545,g21562);
	not 	XG11581 	(g22865,g20330);
	not 	XG11582 	(g22985,g20330);
	not 	XG11583 	(g23011,g20330);
	not 	XG11584 	(g23302,g20330);
	not 	XG11585 	(g23282,g20330);
	not 	XG11586 	(g22995,g20330);
	not 	XG11587 	(g22840,g20330);
	not 	XG11588 	(g23066,g20330);
	not 	XG11589 	(g22974,g20330);
	not 	XG11590 	(g22922,g20330);
	not 	XG11591 	(g22854,g20330);
	not 	XG11592 	(g22866,g20330);
	not 	XG11593 	(g22986,g20330);
	not 	XG11594 	(g23012,g20330);
	not 	XG11595 	(g23406,g20330);
	not 	XG11596 	(g22996,g20330);
	not 	XG11597 	(g23013,g20330);
	not 	XG11598 	(g22903,g20330);
	not 	XG11599 	(g22758,g20330);
	not 	XG11600 	(g22973,g20330);
	not 	XG11601 	(g23245,g20785);
	not 	XG11602 	(g23350,g20785);
	not 	XG11603 	(g23303,g20785);
	not 	XG11604 	(g23283,g20785);
	not 	XG11605 	(g23537,g20785);
	not 	XG11606 	(g23236,g20785);
	not 	XG11607 	(g23222,g20785);
	not 	XG11608 	(g23334,g20785);
	not 	XG11609 	(g23486,g20785);
	not 	XG11610 	(g23256,g20785);
	not 	XG11611 	(g23196,g20785);
	not 	XG11612 	(g23246,g20785);
	not 	XG11613 	(g23473,g20785);
	not 	XG11614 	(g23221,g20785);
	not 	XG11615 	(g23332,g20785);
	not 	XG11616 	(g23515,g20785);
	not 	XG11617 	(g23235,g20785);
	not 	XG11618 	(g23214,g20785);
	not 	XG11619 	(g23333,g20785);
	not 	XG11620 	(g23304,g20785);
	not 	XG11621 	(g23284,g20785);
	not 	XG11622 	(g23215,g20785);
	not 	XG11623 	(g23485,g20785);
	not 	XG11624 	(g23270,g20785);
	not 	XG11625 	(g23271,g20785);
	not 	XG11626 	(g23499,g20785);
	not 	XG11627 	(g23925,g21514);
	not 	XG11628 	(g23505,g21514);
	not 	XG11629 	(g23522,g21514);
	not 	XG11630 	(g23409,g21514);
	not 	XG11631 	(g23905,g21514);
	not 	XG11632 	(g23542,g21514);
	not 	XG11633 	(g23523,g21514);
	not 	XG11634 	(g23543,g21514);
	not 	XG11635 	(g23478,g21514);
	not 	XG11636 	(g23431,g21514);
	not 	XG11637 	(g23456,g21514);
	not 	XG11638 	(g23490,g21514);
	not 	XG11639 	(g23420,g21514);
	not 	XG11640 	(g23629,g21514);
	not 	XG11641 	(g23491,g21514);
	not 	XG11642 	(g23506,g21514);
	not 	XG11643 	(g23541,g21514);
	not 	XG11644 	(g24003,g21514);
	not 	XG11645 	(g23399,g21514);
	not 	XG11646 	(g23432,g21514);
	not 	XG11647 	(g23793,g19074);
	not 	XG11648 	(g23961,g19074);
	not 	XG11649 	(g23769,g19074);
	not 	XG11650 	(g23840,g19074);
	not 	XG11651 	(g22148,g19074);
	not 	XG11652 	(g23841,g19074);
	not 	XG11653 	(g23814,g19074);
	not 	XG11654 	(g23815,g19074);
	not 	XG11655 	(g23876,g19074);
	not 	XG11656 	(g23894,g19074);
	not 	XG11657 	(g23860,g19074);
	not 	XG11658 	(g23859,g19074);
	not 	XG11659 	(g23926,g19074);
	not 	XG11660 	(g22197,g19074);
	not 	XG11661 	(g23927,g19074);
	not 	XG11662 	(g23940,g19074);
	not 	XG11663 	(g23906,g19074);
	not 	XG11664 	(g23941,g19074);
	not 	XG11665 	(g23907,g19074);
	not 	XG11666 	(g23939,g19074);
	not 	XG11667 	(g23893,g19074);
	not 	XG11668 	(g22154,g19074);
	not 	XG11669 	(g23792,g19074);
	not 	XG11670 	(g22177,g19074);
	not 	XG11671 	(g22167,g19074);
	not 	XG11672 	(g22155,g19074);
	not 	XG11673 	(g22201,g19277);
	not 	XG11674 	(g23995,g19277);
	not 	XG11675 	(g22224,g19277);
	not 	XG11676 	(g23881,g19277);
	not 	XG11677 	(g23952,g19277);
	not 	XG11678 	(g23953,g19277);
	not 	XG11679 	(g22303,g19277);
	not 	XG11680 	(g23937,g19277);
	not 	XG11681 	(g23993,g19277);
	not 	XG11682 	(g23916,g19277);
	not 	XG11683 	(g23969,g19277);
	not 	XG11684 	(g23987,g19277);
	not 	XG11685 	(g23898,g19277);
	not 	XG11686 	(g23899,g19277);
	not 	XG11687 	(g22181,g19277);
	not 	XG11688 	(g23849,g19277);
	not 	XG11689 	(g23882,g19277);
	not 	XG11690 	(g23915,g19277);
	not 	XG11691 	(g22200,g19277);
	not 	XG11692 	(g24000,g19277);
	not 	XG11693 	(g22215,g19277);
	not 	XG11694 	(g23994,g19277);
	not 	XG11695 	(g23970,g19277);
	not 	XG11696 	(g23868,g19277);
	not 	XG11697 	(g23869,g19277);
	not 	XG11698 	(g23988,g19277);
	not 	XG11699 	(g23548,g18833);
	not 	XG11700 	(g23549,g18833);
	not 	XG11701 	(g23449,g18833);
	not 	XG11702 	(g23647,g18833);
	not 	XG11703 	(g23482,g18833);
	not 	XG11704 	(g23483,g18833);
	not 	XG11705 	(g23510,g18833);
	not 	XG11706 	(g23986,g18833);
	not 	XG11707 	(g23968,g18833);
	not 	XG11708 	(g24017,g18833);
	not 	XG11709 	(g23648,g18833);
	not 	XG11710 	(g23649,g18833);
	not 	XG11711 	(g23435,g18833);
	not 	XG11712 	(g23732,g18833);
	not 	XG11713 	(g23570,g18833);
	not 	XG11714 	(g23610,g18833);
	not 	XG11715 	(g23571,g18833);
	not 	XG11716 	(g23528,g18833);
	not 	XG11717 	(g23461,g18833);
	not 	XG11718 	(g23611,g18833);
	and 	XG11719 	(g24408,g18946,g23989);
	and 	XG11720 	(g26844,g21418,g25261);
	and 	XG11721 	(g25979,g19650,g24517);
	or 	XG11722 	(g24374,g24004,g19345);
	nand 	XG11723 	(I21978,I21976,g19620);
	nand 	XG11724 	(I22946,I22944,g19620);
	nand 	XG11725 	(I21994,I21992,g19638);
	nand 	XG11726 	(I22974,I22972,g19638);
	or 	XG11727 	(g24276,g18646,g23083);
	or 	XG11728 	(g24277,g18647,g23188);
	or 	XG11729 	(g25613,g18140,g25181);
	or 	XG11730 	(g25603,g18114,g24698);
	or 	XG11731 	(g25604,g18115,g24717);
	or 	XG11732 	(g25607,g18118,g24773);
	or 	XG11733 	(g25606,g18117,g24761);
	or 	XG11734 	(g25736,g18785,g25536);
	nand 	XG11735 	(I22710,g21434,g11915);
	or 	XG11736 	(g24345,g18788,g23606);
	or 	XG11737 	(g24214,g18195,g23471);
	or 	XG11738 	(g24216,g18197,g23416);
	or 	XG11739 	(g25669,g18624,g24657);
	or 	XG11740 	(g25668,g18623,g24646);
	and 	XG11741 	(g26127,g25119,g2236);
	or 	XG11742 	(g24273,g18630,g23166);
	or 	XG11743 	(g24334,g18676,g23991);
	or 	XG11744 	(g24209,g18122,g23415);
	or 	XG11745 	(g24349,g18805,g23646);
	or 	XG11746 	(g24253,g18300,g22525);
	or 	XG11747 	(g24252,g18299,g22518);
	or 	XG11748 	(g24352,g18821,g22157);
	or 	XG11749 	(g25636,g18305,g24507);
	not 	XG11750 	(g21175,I20951);
	or 	XG11751 	(g24348,g18804,g22149);
	or 	XG11752 	(I22267,g20111,g20133,g20236);
	or 	XG11753 	(g24344,g18787,g22145);
	or 	XG11754 	(g25684,g18643,g24983);
	or 	XG11755 	(g26895,g18148,g26783);
	or 	XG11756 	(g24246,g18257,g23372);
	or 	XG11757 	(g24244,g18255,g23349);
	or 	XG11758 	(g25621,g18205,g24523);
	or 	XG11759 	(g24210,g18125,g22900);
	or 	XG11760 	(g24235,g18238,g22632);
	and 	XG11761 	(g25926,g24839,g25005);
	and 	XG11762 	(g25928,g23436,g25022);
	or 	XG11763 	(g25619,g18193,g24961);
	or 	XG11764 	(g24340,g18770,g24016);
	or 	XG11765 	(g25656,g18609,g24945);
	not 	XG11766 	(I21002,g16709);
	not 	XG11767 	(I20999,g16709);
	or 	XG11768 	(g24265,g18560,g22316);
	not 	XG11769 	(I20985,g16300);
	not 	XG11770 	(I20982,g16300);
	or 	XG11771 	(g25627,g18247,g24503);
	or 	XG11772 	(g25750,g18802,g25543);
	or 	XG11773 	(g26917,g18233,g26122);
	or 	XG11774 	(g24433,g22400,g10878);
	or 	XG11775 	(g24337,g18754,g23540);
	or 	XG11776 	(g24338,g18755,g23658);
	not 	XG11777 	(I21019,g17325);
	or 	XG11778 	(g24258,g18311,g22851);
	or 	XG11779 	(g24251,g18296,g22637);
	or 	XG11780 	(g24250,g18295,g22633);
	or 	XG11781 	(g26924,g18291,g26153);
	or 	XG11782 	(g24259,g18312,g23008);
	or 	XG11783 	(g24255,g18308,g22835);
	nand 	XG11784 	(I22892,g21228,g12189);
	or 	XG11785 	(g24239,g18250,g22752);
	or 	XG11786 	(g24335,g18678,g22165);
	nand 	XG11787 	(I22965,g21228,g12288);
	or 	XG11788 	(g26922,g18288,g25902);
	or 	XG11789 	(g24271,g18628,g23451);
	or 	XG11790 	(g24353,g18822,g23682);
	or 	XG11791 	(g24354,g18823,g23775);
	nand 	XG11792 	(I21993,I21992,g7670);
	or 	XG11793 	(g24282,g18657,g23407);
	or 	XG11794 	(g24281,g18656,g23397);
	or 	XG11795 	(g24237,g18242,g22515);
	or 	XG11796 	(g24249,g18294,g22624);
	or 	XG11797 	(g25734,g18782,g25058);
	or 	XG11798 	(g25655,g18607,g24645);
	or 	XG11799 	(g24270,g18614,g23165);
	and 	XG11800 	(g26288,g25309,g2259);
	or 	XG11801 	(g24206,g18110,g23386);
	or 	XG11802 	(g24205,g18109,g23006);
	or 	XG11803 	(g24351,g18807,g23774);
	or 	XG11804 	(g26914,g18227,g25949);
	not 	XG11805 	(g22150,g21280);
	and 	XG11806 	(g26273,g25389,g2122);
	or 	XG11807 	(g25682,g18640,g24658);
	or 	XG11808 	(g25748,g18799,g25078);
	or 	XG11809 	(g25749,g18800,g25094);
	or 	XG11810 	(g25625,g18226,g24553);
	not 	XG11811 	(g19699,I20116);
	and 	XG11812 	(I24704,g24063,g24062,g24061,g21193);
	or 	XG11813 	(g24272,g18629,g23056);
	or 	XG11814 	(g25600,g18111,g24650);
	or 	XG11815 	(g25601,g18112,g24660);
	or 	XG11816 	(g26915,g18230,g25900);
	or 	XG11817 	(g24444,g22400,g10890);
	nand 	XG11818 	(I22899,g21228,g12193);
	and 	XG11819 	(g26158,g25432,g2255);
	not 	XG11820 	(I22211,g21463);
	or 	XG11821 	(g24275,g18645,g23474);
	or 	XG11822 	(g25721,g18766,g25057);
	or 	XG11823 	(g24204,g18108,g22990);
	or 	XG11824 	(g25635,g18293,g24504);
	or 	XG11825 	(g24248,g18286,g22710);
	or 	XG11826 	(g25763,g18817,g25113);
	or 	XG11827 	(g24243,g18254,g22992);
	or 	XG11828 	(g24245,g18256,g22849);
	or 	XG11829 	(g25654,g18606,g24634);
	or 	XG11830 	(g24242,g18253,g22834);
	not 	XG11831 	(I20867,g16216);
	not 	XG11832 	(I20870,g16216);
	or 	XG11833 	(g25628,g18249,g24600);
	or 	XG11834 	(g24260,g18313,g23373);
	or 	XG11835 	(g25638,g18316,g24977);
	or 	XG11836 	(g24262,g18315,g23387);
	or 	XG11837 	(g25720,g18765,g25042);
	or 	XG11838 	(g25747,g18795,g25130);
	or 	XG11839 	(g24460,g22450,g10967);
	nand 	XG11840 	(g24926,g13995,g23357,g20163,g20172);
	and 	XG11841 	(g25580,g24149,g19268);
	or 	XG11842 	(g24278,g18648,g23201);
	or 	XG11843 	(g26923,g18290,g25923);
	or 	XG11844 	(g25608,g18120,g24643);
	or 	XG11845 	(g25612,g18132,g24941);
	or 	XG11846 	(g24266,g18561,g22329);
	or 	XG11847 	(g25639,g18530,g25122);
	not 	XG11848 	(g20695,I20781);
	or 	XG11849 	(g24261,g18314,g22862);
	not 	XG11850 	(I21033,g17221);
	not 	XG11851 	(I21036,g17221);
	not 	XG11852 	(g19458,I19927);
	or 	XG11853 	(g24267,g18611,g23439);
	nand 	XG11854 	(I22822,g21434,g11978);
	nand 	XG11855 	(I21977,I21976,g7680);
	or 	XG11856 	(g24208,g18121,g23404);
	or 	XG11857 	(g24207,g18119,g23396);
	or 	XG11858 	(g25617,g18189,g25466);
	or 	XG11859 	(g25618,g18192,g25491);
	or 	XG11860 	(g25605,g18116,g24743);
	or 	XG11861 	(g24269,g18613,g23131);
	or 	XG11862 	(g24268,g18612,g23025);
	or 	XG11863 	(g24200,g18103,g22831);
	or 	XG11864 	(g24203,g18107,g22982);
	or 	XG11865 	(g24347,g18790,g23754);
	and 	XG11866 	(g26101,g25098,g1760);
	and 	XG11867 	(g26233,g25309,g2279);
	or 	XG11868 	(g25670,g18626,g24967);
	or 	XG11869 	(g24236,g18241,g22489);
	or 	XG11870 	(g24336,g18753,g24012);
	not 	XG11871 	(g18940,I19719);
	or 	XG11872 	(g24233,g18236,g22590);
	or 	XG11873 	(g24234,g18237,g22622);
	or 	XG11874 	(g25667,g18619,g24682);
	or 	XG11875 	(g24471,g22450,g10999);
	or 	XG11876 	(g24211,g18138,g23572);
	or 	XG11877 	(g24341,g18771,g23564);
	or 	XG11878 	(g24342,g18772,g23691);
	or 	XG11879 	(g24232,g18228,g22686);
	or 	XG11880 	(g24201,g18104,g22848);
	or 	XG11881 	(g25602,g18113,g24673);
	or 	XG11882 	(g25634,g18284,g24559);
	nand 	XG11883 	(I22753,g21434,g11937);
	and 	XG11884 	(g25922,g20065,g24959);
	and 	XG11885 	(g25924,g16846,g24976);
	or 	XG11886 	(g25611,g18128,g24931);
	or 	XG11887 	(g25764,g18819,g25551);
	nand 	XG11888 	(I22683,g21434,g11893);
	or 	XG11889 	(g25722,g18768,g25530);
	not 	XG11890 	(I20819,g17088);
	not 	XG11891 	(I20816,g17088);
	or 	XG11892 	(g24215,g18196,g23484);
	or 	XG11893 	(g24799,g23921,g23901);
	or 	XG11894 	(g25733,g18778,g25108);
	and 	XG11895 	(I27528,g24120,g24119,g24118,g20998);
	and 	XG11896 	(I24709,g24070,g24069,g24068,g21256);
	or 	XG11897 	(g24346,g18789,g23725);
	or 	XG11898 	(g25681,g18636,g24710);
	not 	XG11899 	(I22009,g21269);
	not 	XG11900 	(g23191,I22289);
	not 	XG11901 	(I23324,g21697);
	not 	XG11902 	(I23303,g21669);
	not 	XG11903 	(I23312,g21681);
	not 	XG11904 	(I23318,g21689);
	not 	XG11905 	(I23300,g21665);
	not 	XG11906 	(I23315,g21685);
	not 	XG11907 	(I23306,g21673);
	not 	XG11908 	(I23309,g21677);
	not 	XG11909 	(I23321,g21693);
	or 	XG11910 	(g25761,g18812,g25152);
	or 	XG11911 	(g24578,g23825,g2882);
	or 	XG11912 	(g24782,g23872,g23857);
	or 	XG11913 	(g24447,g22450,g10948);
	and 	XG11914 	(I24679,g24028,g24027,g24026,g19968);
	or 	XG11915 	(g25610,g18127,g24923);
	or 	XG11916 	(g25708,g18751,g25526);
	not 	XG11917 	(I20233,g17487);
	or 	XG11918 	(g24263,g18529,g23497);
	nor 	XG11919 	(g24575,g23514,g23498);
	and 	XG11920 	(g26272,g25470,g2036);
	not 	XG11921 	(g18926,I19707);
	or 	XG11922 	(g25609,g18126,g24915);
	or 	XG11923 	(g25630,g18263,g24532);
	or 	XG11924 	(g24247,g18259,g22623);
	or 	XG11925 	(g25719,g18761,g25089);
	or 	XG11926 	(g24231,g18201,g22589);
	nand 	XG11927 	(I22799,g21434,g11960);
	and 	XG11928 	(g26310,g25389,g2102);
	and 	XG11929 	(g25965,g24980,g2208);
	nor 	XG11930 	(g24497,g23553,g23533);
	or 	XG11931 	(g25615,g18162,g24803);
	or 	XG11932 	(g26916,g18232,g25916);
	not 	XG11933 	(I19671,g15932);
	not 	XG11934 	(I19674,g15932);
	nand 	XG11935 	(I22945,I22944,g9492);
	and 	XG11936 	(g26205,g25492,g2098);
	and 	XG11937 	(g26230,g25385,g1768);
	or 	XG11938 	(g26921,g18285,g25955);
	not 	XG11939 	(g26615,g25432);
	not 	XG11940 	(g26702,g25309);
	not 	XG11941 	(g26682,g25309);
	not 	XG11942 	(g26765,g25309);
	not 	XG11943 	(g21366,I21100);
	nand 	XG11944 	(I22792,g21434,g11956);
	or 	XG11945 	(g24350,g18806,g23755);
	not 	XG11946 	(I20753,g16677);
	not 	XG11947 	(I20750,g16677);
	not 	XG11948 	(g26679,g25385);
	not 	XG11949 	(g19720,I20130);
	not 	XG11950 	(I20861,g16960);
	not 	XG11951 	(I20864,g16960);
	or 	XG11952 	(g24457,g22400,g10902);
	nand 	XG11953 	(I22717,g21434,g11916);
	or 	XG11954 	(g25629,g18258,g24962);
	not 	XG11955 	(I20957,g16228);
	not 	XG11956 	(I20954,g16228);
	not 	XG11957 	(g26655,g25492);
	not 	XG11958 	(g26803,g25389);
	not 	XG11959 	(g26758,g25389);
	not 	XG11960 	(g26732,g25389);
	not 	XG11961 	(I20650,g17010);
	not 	XG11962 	(I20647,g17010);
	or 	XG11963 	(g24202,g18106,g22899);
	or 	XG11964 	(g25705,g18744,g25069);
	not 	XG11965 	(I22124,g21300);
	or 	XG11966 	(g24355,g18824,g23799);
	or 	XG11967 	(g25626,g18235,g24499);
	or 	XG11968 	(g24468,g22400,g10925);
	or 	XG11969 	(g25835,g23855,g25367);
	or 	XG11970 	(g25762,g18816,g25095);
	and 	XG11971 	(g25579,g24147,g19422);
	or 	XG11972 	(g24343,g18773,g23724);
	or 	XG11973 	(g25867,g23884,g25449);
	or 	XG11974 	(g25735,g18783,g25077);
	or 	XG11975 	(g25706,g18748,g25030);
	or 	XG11976 	(g24274,g18631,g23187);
	not 	XG11977 	(I21831,g19127);
	not 	XG11978 	(I22470,g21326);
	not 	XG11979 	(I22589,g21340);
	not 	XG11980 	(I22240,g20086);
	not 	XG11981 	(I22275,g20127);
	not 	XG11982 	(I22264,g20100);
	not 	XG11983 	(g26731,g25470);
	nand 	XG11984 	(g24574,g22687,g22709);
	nand 	XG11985 	(g24591,g22642,g22833);
	or 	XG11986 	(g25906,g24014,g25559);
	or 	XG11987 	(g25683,g18641,g24669);
	or 	XG11988 	(g25707,g18749,g25041);
	not 	XG11989 	(I20747,g17141);
	not 	XG11990 	(I20744,g17141);
	or 	XG11991 	(g25637,g18307,g24618);
	or 	XG11992 	(g25653,g18602,g24664);
	or 	XG11993 	(g24339,g18756,g23690);
	not 	XG11994 	(I20321,g16920);
	not 	XG11995 	(I20318,g16920);
	and 	XG11996 	(g23708,g9104,g19050);
	and 	XG11997 	(g23599,g9104,g19050);
	and 	XG11998 	(g23675,g9104,g19050);
	and 	XG11999 	(g23828,g19128,g9104);
	and 	XG12000 	(g23121,g9104,g19128);
	and 	XG12001 	(g22689,g9104,g18918);
	and 	XG12002 	(g22876,g9104,g20136);
	and 	XG12003 	(g22942,g20219,g9104);
	and 	XG12004 	(g22670,g9104,g20114);
	and 	XG12005 	(g23314,g19200,g9104);
	and 	XG12006 	(g23076,g9104,g19128);
	and 	XG12007 	(g23639,g9104,g19050);
	and 	XG12008 	(g23293,g19200,g9104);
	and 	XG12009 	(g23148,g9104,g19128);
	and 	XG12010 	(g23958,g19200,g9104);
	and 	XG12011 	(g23742,g9104,g19128);
	and 	XG12012 	(g23802,g19050,g9104);
	nand 	XG12013 	(g22885,g20154,g9104);
	nand 	XG12014 	(g22908,g20175,g9104);
	and 	XG12015 	(g26229,g25275,g1724);
	nand 	XG12016 	(g22941,g2970,g20219);
	and 	XG12017 	(g26311,g25400,g2527);
	not 	XG12018 	(I21930,g21297);
	not 	XG12019 	(I22302,g19353);
	not 	XG12020 	(I21911,g21278);
	not 	XG12021 	(I22316,g19361);
	not 	XG12022 	(I22327,g19367);
	not 	XG12023 	(I22353,g19375);
	not 	XG12024 	(I21918,g21290);
	not 	XG12025 	(I22343,g19371);
	and 	XG12026 	(g25970,g24991,g1792);
	and 	XG12027 	(g26251,g25341,g1988);
	and 	XG12028 	(g26324,g25439,g2661);
	nand 	XG12029 	(g23266,g2894,g18918);
	and 	XG12030 	(g25959,g24963,g1648);
	nand 	XG12031 	(I22844,g21228,g12113);
	or 	XG12032 	(g22516,g12817,g21559);
	nand 	XG12033 	(g22668,g2912,g20219);
	and 	XG12034 	(g26160,g25138,g2453);
	and 	XG12035 	(g26104,g25101,g2250);
	or 	XG12036 	(g24478,g22450,g11003);
	and 	XG12037 	(g26177,g25154,g2079);
	nand 	XG12038 	(g22661,g94,g20136);
	and 	XG12039 	(g25991,g25023,g2060);
	nand 	XG12040 	(g22853,g2922,g20219);
	nand 	XG12041 	(g22688,g2936,g20219);
	and 	XG12042 	(g26091,g25082,g1691);
	and 	XG12043 	(g26254,g25349,g2413);
	and 	XG12044 	(g26291,g25439,g2681);
	and 	XG12045 	(g25957,g24960,g17190);
	nand 	XG12046 	(g22715,g2999,g20114);
	and 	XG12047 	(g26285,g25300,g1834);
	and 	XG12048 	(g26253,g25435,g2327);
	and 	XG12049 	(g25981,g25007,g2051);
	nand 	XG12050 	(I22929,g21228,g12223);
	nand 	XG12051 	(I22760,g21434,g11939);
	or 	XG12052 	(g25836,g23856,g25368);
	or 	XG12053 	(g25877,g23919,g25502);
	and 	XG12054 	(g26204,g25275,g1720);
	and 	XG12055 	(g26176,g25467,g1964);
	and 	XG12056 	(g26286,g25389,g2126);
	not 	XG12057 	(g26820,I25534);
	and 	XG12058 	(g26250,g25429,g1902);
	nand 	XG12059 	(g22852,g2856,g18957);
	nand 	XG12060 	(g22713,g2890,g20114);
	and 	XG12061 	(g26124,g25116,g1811);
	and 	XG12062 	(g26249,g25300,g1858);
	or 	XG12063 	(g25819,g23836,g25323);
	nand 	XG12064 	(g22921,g2950,g20219);
	and 	XG12065 	(g26303,g25439,g2685);
	and 	XG12066 	(g26157,g25136,g2093);
	nand 	XG12067 	(g22757,g7891,g20114);
	and 	XG12068 	(g25972,g24993,g2217);
	and 	XG12069 	(g26207,g25170,g2638);
	and 	XG12070 	(g26156,g25135,g2028);
	and 	XG12071 	(g26100,g25097,g1677);
	and 	XG12072 	(g26090,g25081,g1624);
	and 	XG12073 	(g26154,g25426,g1830);
	and 	XG12074 	(g26341,g20105,g24746);
	and 	XG12075 	(g24554,g19541,g22490);
	and 	XG12076 	(g25964,g24979,g1783);
	nand 	XG12077 	(I22864,g21228,g12146);
	nand 	XG12078 	(g22984,g2868,g20114);
	and 	XG12079 	(g26252,g25309,g2283);
	and 	XG12080 	(g26845,g21426,g24391);
	and 	XG12081 	(g26684,g20673,g25407);
	and 	XG12082 	(g26713,g20714,g25447);
	and 	XG12083 	(g26711,g20713,g25446);
	and 	XG12084 	(g26635,g20617,g25321);
	and 	XG12085 	(g25951,g19565,g24500);
	nand 	XG12086 	(g23195,g37,g20136);
	and 	XG12087 	(g26103,g25100,g2185);
	nand 	XG12088 	(I20188,I20187,g16272);
	nand 	XG12089 	(I20222,I20221,g16272);
	and 	XG12090 	(g26179,g25155,g2504);
	and 	XG12091 	(g26611,g20580,g24935);
	or 	XG12092 	(g22487,g12794,g21512);
	and 	XG12093 	(g26102,g25099,g1825);
	and 	XG12094 	(g25946,g19537,g24496);
	and 	XG12095 	(g26178,g25473,g2389);
	and 	XG12096 	(g25925,g23234,g24990);
	and 	XG12097 	(g25927,g20375,g25004);
	and 	XG12098 	(g24797,g19960,g22872);
	nor 	XG12099 	(g24514,g23657,g23619);
	nor 	XG12100 	(g24508,g23618,g23577);
	nor 	XG12101 	(g24494,g23532,g23513);
	not 	XG12102 	(g26681,g25396);
	nand 	XG12103 	(I22871,g21228,g12150);
	and 	XG12104 	(g26231,g25300,g1854);
	nand 	XG12105 	(g22651,g2873,g20114);
	and 	XG12106 	(g25904,g24791,g14001);
	and 	XG12107 	(g26387,g20231,g24813);
	and 	XG12108 	(g27160,g26340,g14163);
	and 	XG12109 	(g24997,g10419,g22929);
	and 	XG12110 	(g25026,g10503,g22929);
	and 	XG12111 	(g24984,g12818,g22929);
	nand 	XG12112 	(g24890,g22929,g13852);
	nand 	XG12113 	(g24936,g14029,g23379,g20173,g20186);
	nor 	XG12114 	(g24619,g23581,g23554);
	and 	XG12115 	(g27268,g19733,g25942);
	and 	XG12116 	(g26289,g25400,g2551);
	or 	XG12117 	(g24841,g23998,g21420);
	and 	XG12118 	(g26799,g21068,g25247);
	not 	XG12119 	(g26720,g25275);
	not 	XG12120 	(g26654,g25275);
	not 	XG12121 	(g26672,g25275);
	not 	XG12122 	(I22149,g21036);
	not 	XG12123 	(g26743,g25476);
	nand 	XG12124 	(I22936,g21228,g12226);
	and 	XG12125 	(g27255,g19689,g25936);
	nand 	XG12126 	(g22712,g2864,g18957);
	and 	XG12127 	(g26778,g20923,g25501);
	nand 	XG12128 	(g23210,g2882,g18957);
	nand 	XG12129 	(g22666,g2878,g18957);
	and 	XG12130 	(g27249,g19678,g25929);
	nand 	XG12131 	(g22839,g2988,g20114);
	not 	XG12132 	(g26631,g25467);
	and 	XG12133 	(g27263,g19713,g25940);
	nand 	XG12134 	(I20166,I20165,g16246);
	nand 	XG12135 	(I20204,I20203,g16246);
	or 	XG12136 	(g27456,g24607,g25978);
	and 	XG12137 	(g23254,g20110,g20056);
	not 	XG12138 	(I24558,g23777);
	not 	XG12139 	(g26683,g25514);
	nand 	XG12140 	(g22940,g2860,g18918);
	not 	XG12141 	(g27242,g26183);
	or 	XG12142 	(g24853,g24001,g21452);
	or 	XG12143 	(g24821,g23990,g21404);
	or 	XG12144 	(g24840,g23996,g21419);
	or 	XG12145 	(g24907,g24015,g21558);
	and 	XG12146 	(g27269,g19734,g25943);
	and 	XG12147 	(g26302,g25349,g2393);
	not 	XG12148 	(g26777,g25439);
	not 	XG12149 	(g26812,g25439);
	not 	XG12150 	(g26792,g25439);
	not 	XG12151 	(g26754,g25300);
	not 	XG12152 	(g26693,g25300);
	not 	XG12153 	(g26680,g25300);
	not 	XG12154 	(g26614,g25426);
	nor 	XG12155 	(g23956,g20114,g20136,g18918,g18957);
	not 	XG12156 	(I21941,g18918);
	nor 	XG12157 	(g22405,g20114,g20136,g18957);
	not 	XG12158 	(g22994,g20436);
	not 	XG12159 	(g22756,g20436);
	not 	XG12160 	(g22714,g20436);
	not 	XG12161 	(I22143,g20189);
	and 	XG12162 	(g26808,g21185,g25521);
	and 	XG12163 	(g26271,g25341,g1992);
	and 	XG12164 	(g27378,g20052,g26089);
	and 	XG12165 	(g26275,g25349,g2417);
	and 	XG12166 	(g26290,g25498,g2595);
	nand 	XG12167 	(I22973,I22972,g9657);
	nand 	XG12168 	(g23010,g2984,g20516);
	nand 	XG12169 	(I20189,I20187,g1333);
	or 	XG12170 	(I22880,g21351,g21356,g21509);
	not 	XG12171 	(g26710,g25349);
	not 	XG12172 	(g26788,g25349);
	not 	XG12173 	(g26736,g25349);
	not 	XG12174 	(g26632,g25473);
	nand 	XG12175 	(g14677,I16780,I16779);
	and 	XG12176 	(g23265,g20132,g20069);
	or 	XG12177 	(I22280,g20134,g20150,g20271);
	or 	XG12178 	(I22830,g21307,g21338,g21429);
	nand 	XG12179 	(g22643,g18954,g20136);
	nand 	XG12180 	(g22755,g18984,g20136);
	nand 	XG12181 	(g22754,g19376,g20114);
	not 	XG12182 	(I21838,g19263);
	or 	XG12183 	(I22852,g21339,g21350,g21459);
	or 	XG12184 	(g25885,g23957,g25522);
	nand 	XG12185 	(I20223,I20221,g11170);
	not 	XG12186 	(g25766,g24439);
	not 	XG12187 	(g26709,g25435);
	and 	XG12188 	(g24546,g19523,g22447);
	or 	XG12189 	(g25878,g23920,g25503);
	or 	XG12190 	(g25868,g23885,g25450);
	and 	XG12191 	(g27254,g19688,g25935);
	and 	XG12192 	(g27275,g19745,g25945);
	not 	XG12193 	(g26776,g25498);
	not 	XG12194 	(g26700,g25429);
	not 	XG12195 	(g26769,g25400);
	not 	XG12196 	(g26804,g25400);
	not 	XG12197 	(g26744,g25400);
	and 	XG12198 	(g27264,g19714,g25941);
	not 	XG12199 	(g26784,g25341);
	not 	XG12200 	(g26701,g25341);
	not 	XG12201 	(g26724,g25341);
	and 	XG12202 	(g24817,g7235,g22929);
	and 	XG12203 	(g24420,g18980,g23997);
	or 	XG12204 	(I22912,g21357,g21364,g21555);
	and 	XG12205 	(g23218,g16530,g20200);
	and 	XG12206 	(g26277,g25400,g2547);
	nand 	XG12207 	(g22837,g2907,g20219);
	and 	XG12208 	(g26300,g25341,g1968);
	and 	XG12209 	(g26234,g25514,g2657);
	nand 	XG12210 	(g22874,g2844,g18918);
	nor 	XG12211 	(g26338,g24825,g8458);
	and 	XG12212 	(g25980,g25006,g1926);
	nor 	XG12213 	(g26309,g24825,g8575);
	or 	XG12214 	(g27533,g24659,g26078);
	and 	XG12215 	(g25992,g25024,g2485);
	and 	XG12216 	(g26203,g25337,g1632);
	and 	XG12217 	(g25971,g24992,g1917);
	nand 	XG12218 	(g26352,g11679,g24875,g744);
	and 	XG12219 	(g25909,g24875,g8745);
	and 	XG12220 	(g25993,g25025,g2610);
	nand 	XG12221 	(g22875,g2980,g20516);
	and 	XG12222 	(g27820,g25932,g7670);
	or 	XG12223 	(g25545,g20658,g23551);
	or 	XG12224 	(g27484,g24628,g25988);
	nand 	XG12225 	(g23281,g2898,g18957);
	nand 	XG12226 	(g22836,g2852,g18918);
	not 	XG12227 	(g25930,I25028);
	nand 	XG12228 	(g22638,g2886,g18957);
	nand 	XG12229 	(g25888,g24439,g914);
	and 	XG12230 	(g26572,g24439,g7443);
	and 	XG12231 	(g25973,g24994,g2342);
	and 	XG12232 	(g26514,g25564,g7400);
	nand 	XG12233 	(g22838,g2960,g20219);
	nor 	XG12234 	(g26267,g24732,g8033);
	or 	XG12235 	(I22298,g20151,g20161,g20371);
	or 	XG12236 	(g27233,g24451,g25876);
	nor 	XG12237 	(g26298,g24825,g8297);
	or 	XG12238 	(g27566,g24713,g26119);
	nand 	XG12239 	(g22902,g2848,g18957);
	and 	XG12240 	(g26128,g25120,g2319);
	and 	XG12241 	(g26159,g25137,g2370);
	nor 	XG12242 	(g26247,g24732,g7995);
	and 	XG12243 	(g26276,g25476,g2461);
	and 	XG12244 	(g26544,g24357,g7446);
	or 	XG12245 	(g27575,g24731,g26147);
	and 	XG12246 	(g27965,g13117,g25834);
	not 	XG12247 	(I25750,g26823);
	or 	XG12248 	(g27243,g24475,g25884);
	and 	XG12249 	(g26270,g25275,g1700);
	not 	XG12250 	(g24964,I24128);
	and 	XG12251 	(g26051,g14169,g24896);
	or 	XG12252 	(g27543,g24670,g26085);
	not 	XG12253 	(g27038,g25932);
	nand 	XG12254 	(I20167,I20165,g990);
	nor 	XG12255 	(g26296,g24732,g8287);
	or 	XG12256 	(g27663,g24820,g26323);
	and 	XG12257 	(g26024,g25039,g2619);
	and 	XG12258 	(g26181,g25157,g2652);
	and 	XG12259 	(g26232,g25396,g2193);
	nor 	XG12260 	(g26098,g24732,g9073);
	and 	XG12261 	(g26123,g25382,g1696);
	nand 	XG12262 	(I20205,I20203,g11147);
	and 	XG12263 	(g26180,g25156,g2587);
	or 	XG12264 	(g27556,g24687,g26097);
	nand 	XG12265 	(g27679,g26685,g25186);
	and 	XG12266 	(g25982,g25008,g2351);
	or 	XG12267 	(g27239,g24465,g25881);
	or 	XG12268 	(g27509,g24640,g26023);
	or 	XG12269 	(g27147,g24399,g25802);
	nor 	XG12270 	(g26346,g24825,g8522);
	and 	XG12271 	(g26125,g25117,g1894);
	or 	XG12272 	(g26299,g22665,g24551);
	or 	XG12273 	(g27584,g24758,g26165);
	and 	XG12274 	(g26161,g25139,g2518);
	nor 	XG12275 	(g26297,g24825,g8519);
	and 	XG12276 	(g26155,g25134,g1945);
	and 	XG12277 	(g26126,g25118,g1959);
	not 	XG12278 	(g25222,I24400);
	and 	XG12279 	(g25983,g25009,g2476);
	and 	XG12280 	(g25963,g24978,g1657);
	nor 	XG12281 	(g26268,g24825,g283);
	nor 	XG12282 	(g26330,g24825,g8631);
	and 	XG12283 	(g26129,g25121,g2384);
	and 	XG12284 	(g26206,g25495,g2523);
	or 	XG12285 	(g24879,g24009,g21465);
	or 	XG12286 	(g24919,g22143,g21606);
	or 	XG12287 	(g24854,g24002,g21453);
	not 	XG12288 	(g27565,g26645);
	not 	XG12289 	(g27415,g26382);
	and 	XG12290 	(g25883,g24699,g13728);
	not 	XG12291 	(g26284,g24875);
	not 	XG12292 	(g27592,g26715);
	or 	XG12293 	(g27179,g24409,g25816);
	or 	XG12294 	(g27506,g24639,g26021);
	or 	XG12295 	(g27453,g24606,g25976);
	and 	XG12296 	(g26092,g25083,g9766);
	nor 	XG12297 	(g26609,g24732,g146);
	nor 	XG12298 	(g26598,g24732,g13756,g8990);
	nor 	XG12299 	(g26628,g24732,g8990);
	not 	XG12300 	(g26607,g25382);
	or 	XG12301 	(g25539,g20628,g23531);
	or 	XG12302 	(g25937,g22216,g24406);
	nand 	XG12303 	(g27705,g26782,g25237);
	nand 	XG12304 	(g24583,g22711,g22753);
	nand 	XG12305 	(g24609,g22650,g22850);
	or 	XG12306 	(g27426,g24588,g25967);
	and 	XG12307 	(g24502,g13223,g23428);
	or 	XG12308 	(g27524,g24649,g26050);
	or 	XG12309 	(g27232,g24450,g25874);
	not 	XG12310 	(g26656,g25495);
	nor 	XG12311 	(g26649,g24732,g9037);
	not 	XG12312 	(g26653,g25337);
	nand 	XG12313 	(g27306,g26235,g24787);
	not 	XG12314 	(g24506,I23711);
	or 	XG12315 	(g27133,g24392,g25788);
	or 	XG12316 	(g26512,g23130,g24786);
	or 	XG12317 	(g27226,g24436,g25872);
	not 	XG12318 	(g27554,g26625);
	not 	XG12319 	(g27583,g26686);
	nor 	XG12320 	(g27629,g12259,g26382,g8891);
	and 	XG12321 	(g27145,g26382,g14121);
	or 	XG12322 	(g27544,g24671,g26087);
	or 	XG12323 	(g27487,g24629,g25990);
	or 	XG12324 	(g26361,g22991,g24674);
	or 	XG12325 	(g26386,g23023,g24719);
	or 	XG12326 	(g26392,g23050,g24745);
	or 	XG12327 	(g27403,g24581,g25962);
	or 	XG12328 	(g26359,g22939,g24651);
	or 	XG12329 	(g27555,g24686,g26095);
	or 	XG12330 	(g26377,g23007,g24700);
	or 	XG12331 	(g27429,g24589,g25969);
	not 	XG12332 	(g26634,g25317);
	and 	XG12333 	(g26602,g24453,g7487);
	nand 	XG12334 	(g25895,g24453,g1259);
	or 	XG12335 	(g25910,g22142,g25565);
	or 	XG12336 	(g27567,g24714,g26121);
	or 	XG12337 	(I22958,g21365,g21386,g21603);
	not 	XG12338 	(g27237,g26162);
	or 	XG12339 	(g27238,g24464,g25879);
	or 	XG12340 	(g27182,g24410,g25818);
	and 	XG12341 	(g27020,g25852,g4601);
	or 	XG12342 	(g27150,g24400,g25804);
	or 	XG12343 	(g26396,g23062,g24762);
	or 	XG12344 	(g26422,g23104,g24774);
	nand 	XG12345 	(I23119,I23118,g20076);
	and 	XG12346 	(g27821,g25892,g7680);
	nand 	XG12347 	(g27670,g26666,g25172);
	or 	XG12348 	(g26349,g13409,g24630);
	not 	XG12349 	(g25773,g24453);
	or 	XG12350 	(g27574,g24730,g26145);
	not 	XG12351 	(g27015,g26869);
	or 	XG12352 	(g26972,g25229,g26780);
	or 	XG12353 	(g27205,g24421,g25833);
	nand 	XG12354 	(g27295,g26208,g24776);
	nand 	XG12355 	(g27693,g26752,g25216);
	not 	XG12356 	(g27991,g25852);
	nand 	XG12357 	(I23120,I23118,g417);
	not 	XG12358 	(g27573,g26667);
	nand 	XG12359 	(g27687,g26714,g25200);
	not 	XG12360 	(g27245,g26209);
	nand 	XG12361 	(g27317,g26255,g24793);
	nand 	XG12362 	(g26745,g25317,g6856);
	and 	XG12363 	(g26182,g25317,g9978);
	and 	XG12364 	(g24638,g19690,g22763);
	not 	XG12365 	(g22228,I21810);
	not 	XG12366 	(g22550,I21922);
	and 	XG12367 	(g24627,g19679,g22763);
	not 	XG12368 	(g22722,I22031);
	not 	XG12369 	(g22594,I21934);
	not 	XG12370 	(I23348,g23384);
	not 	XG12371 	(I23378,g23426);
	not 	XG12372 	(g25282,g22763);
	not 	XG12373 	(g25183,g22763);
	not 	XG12374 	(g25283,g22763);
	not 	XG12375 	(g25274,g22763);
	not 	XG12376 	(g25542,g22763);
	not 	XG12377 	(g25208,g22763);
	not 	XG12378 	(g25209,g22763);
	not 	XG12379 	(g24996,g22763);
	not 	XG12380 	(g25193,g22763);
	not 	XG12381 	(g25340,g22763);
	not 	XG12382 	(g24981,g22763);
	not 	XG12383 	(g24770,g22763);
	not 	XG12384 	(g25556,g22763);
	not 	XG12385 	(g25169,g22763);
	not 	XG12386 	(g25557,g22763);
	not 	XG12387 	(g25243,g22763);
	not 	XG12388 	(g25307,g22763);
	not 	XG12389 	(g25550,g22763);
	not 	XG12390 	(g25196,g22763);
	not 	XG12391 	(I24434,g22763);
	not 	XG12392 	(g25211,g22763);
	not 	XG12393 	(g25226,g22763);
	not 	XG12394 	(g25562,g22763);
	not 	XG12395 	(g25227,g22763);
	not 	XG12396 	(g25534,g22763);
	not 	XG12397 	(g25388,g22763);
	not 	XG12398 	(g25262,g22763);
	not 	XG12399 	(g24966,g22763);
	not 	XG12400 	(g25535,g22763);
	not 	XG12401 	(g25541,g22763);
	not 	XG12402 	(g25263,g22763);
	not 	XG12403 	(g25399,g22763);
	not 	XG12404 	(g24995,g22763);
	not 	XG12405 	(g25184,g22763);
	not 	XG12406 	(g25348,g22763);
	not 	XG12407 	(g25438,g22763);
	not 	XG12408 	(g25194,g22763);
	not 	XG12409 	(g24756,g22763);
	not 	XG12410 	(g25195,g22763);
	not 	XG12411 	(g24982,g22763);
	not 	XG12412 	(g25308,g22763);
	not 	XG12413 	(g25224,g22763);
	not 	XG12414 	(g25529,g22763);
	not 	XG12415 	(g25316,g22763);
	not 	XG12416 	(g25299,g22763);
	not 	XG12417 	(g25245,g22763);
	not 	XG12418 	(g25549,g22763);
	not 	XG12419 	(g25011,g22763);
	not 	XG12420 	(g25212,g22763);
	not 	XG12421 	(g25182,g22763);
	not 	XG12422 	(g25356,g22763);
	not 	XG12423 	(I23366,g23321);
	not 	XG12424 	(I23387,g23394);
	not 	XG12425 	(I23360,g23360);
	or 	XG12426 	(g26866,g24363,g20242,g20204);
	not 	XG12427 	(I23327,g22647);
	not 	XG12428 	(I23375,g23403);
	not 	XG12429 	(I23357,g23359);
	not 	XG12430 	(I23333,g22683);
	not 	XG12431 	(I23354,g23277);
	not 	XG12432 	(I23399,g23450);
	not 	XG12433 	(I23336,g22721);
	not 	XG12434 	(I23363,g23385);
	not 	XG12435 	(I23330,g22658);
	not 	XG12436 	(I23381,g23322);
	not 	XG12437 	(I23384,g23362);
	not 	XG12438 	(I23369,g23347);
	not 	XG12439 	(I23393,g23414);
	not 	XG12440 	(g24718,g22182);
	not 	XG12441 	(I23998,g22182);
	not 	XG12442 	(I24008,g22182);
	not 	XG12443 	(I24022,g22182);
	not 	XG12444 	(I24041,g22182);
	nor 	XG12445 	(g25540,g22360,g22409);
	nor 	XG12446 	(g24383,g22360,g22409);
	not 	XG12447 	(I24191,g22360);
	not 	XG12448 	(I24215,g22360);
	not 	XG12449 	(I24078,g22360);
	not 	XG12450 	(I23342,g23299);
	not 	XG12451 	(I23372,g23361);
	not 	XG12452 	(I23396,g23427);
	not 	XG12453 	(I23351,g23263);
	not 	XG12454 	(I23390,g23395);
	not 	XG12455 	(I23339,g23232);
	not 	XG12456 	(I23345,g23320);
	not 	XG12457 	(I24089,g22409);
	not 	XG12458 	(I24228,g22409);
	not 	XG12459 	(I24038,g22202);
	not 	XG12460 	(I24060,g22202);
	not 	XG12461 	(g24744,g22202);
	and 	XG12462 	(g25573,I24705,I24704);
	or 	XG12463 	(I23756,g23511,g23494,g23480,g23457);
	or 	XG12464 	(g26879,g25581,g25580);
	or 	XG12465 	(g24641,g22159,g22151);
	or 	XG12466 	(I26742,g23481,g23458,g23445,g23430);
	and 	XG12467 	(g25574,I24710,I24709);
	or 	XG12468 	(g26363,g24965,g2965);
	and 	XG12469 	(g25568,I24680,I24679);
	or 	XG12470 	(I23755,g23444,g22980,g22927,g22904);
	and 	XG12471 	(g25571,I24695,I24694);
	not 	XG12472 	(I24781,g24264);
	or 	XG12473 	(g26878,g25579,g25578);
	or 	XG12474 	(g24715,g22207,g22189);
	and 	XG12475 	(g25572,I24700,I24699);
	and 	XG12476 	(g25570,I24690,I24689);
	and 	XG12477 	(g25569,I24685,I24684);
	and 	XG12478 	(g25567,I24675,I24674);
	not 	XG12479 	(g20050,I20321);
	or 	XG12480 	(I25736,g20277,g22150,g12);
	nor 	XG12481 	(g22536,g19720,g1379);
	or 	XG12482 	(g24946,g8130,g22409,g22360);
	and 	XG12483 	(g24904,g23279,g11761);
	and 	XG12484 	(g25331,I24508,g22194,g5366);
	or 	XG12485 	(g26721,g24444,g10776);
	or 	XG12486 	(g26785,g24468,g10776);
	or 	XG12487 	(g26766,g24460,g10776);
	or 	XG12488 	(g26755,g24457,g10776);
	or 	XG12489 	(g26789,g24471,g10776);
	or 	XG12490 	(g26733,g24447,g10776);
	or 	XG12491 	(g26690,g24433,g10776);
	and 	XG12492 	(g24794,g23138,g11414);
	and 	XG12493 	(g24777,g23066,g11345);
	and 	XG12494 	(g25187,g23629,g12296);
	and 	XG12495 	(g24729,g23018,g22719);
	and 	XG12496 	(g25201,g23665,g12346);
	and 	XG12497 	(g25091,g23492,g12830);
	not 	XG12498 	(g20653,I20747);
	and 	XG12499 	(g24884,I24051,g23555,g3401);
	and 	XG12500 	(g25045,g23448,g17525);
	and 	XG12501 	(g25462,I24585,g22300,g6404);
	and 	XG12502 	(g27327,g26732,g2116);
	and 	XG12503 	(g27332,g26758,g12538);
	and 	XG12504 	(g24788,g23111,g11384);
	and 	XG12505 	(g24865,g23253,g11323);
	and 	XG12506 	(g27086,g22495,g25836);
	and 	XG12507 	(g27119,g22542,g25877);
	not 	XG12508 	(g23154,I22264);
	not 	XG12509 	(g23172,I22275);
	not 	XG12510 	(g23088,I22240);
	not 	XG12511 	(g23462,I22589);
	not 	XG12512 	(g23363,I22470);
	not 	XG12513 	(g22319,I21831);
	nor 	XG12514 	(g22399,g19720,g1367);
	nor 	XG12515 	(g22537,g1367,g19720);
	and 	XG12516 	(g25104,g23504,g16800);
	and 	XG12517 	(g24864,g22305,g11201);
	and 	XG12518 	(g27097,g22526,g25867);
	and 	XG12519 	(g25179,g23611,g16928);
	nand 	XG12520 	(I22755,I22753,g21434);
	nand 	XG12521 	(I22794,I22792,g21434);
	nand 	XG12522 	(I22719,I22717,g21434);
	nand 	XG12523 	(I22824,I22822,g21434);
	nand 	XG12524 	(I22801,I22799,g21434);
	nand 	XG12525 	(I22685,I22683,g21434);
	nand 	XG12526 	(I22712,I22710,g21434);
	and 	XG12527 	(g24892,g23264,g11559);
	and 	XG12528 	(g24706,g22996,g15910);
	nor 	XG12529 	(g22517,g1345,g19720);
	nor 	XG12530 	(g22523,g19720,g1345);
	and 	XG12531 	(g27083,g22456,g25819);
	nand 	XG12532 	(I23985,g482,g22182);
	and 	XG12533 	(g25059,g23460,g20870);
	and 	XG12534 	(g27085,g22494,g25835);
	not 	XG12535 	(g22923,I22124);
	or 	XG12536 	(g24968,g23389,g22409,g22360);
	and 	XG12537 	(g25173,g23589,g12234);
	and 	XG12538 	(g25238,g23732,g12466);
	or 	XG12539 	(g27571,g24723,g26127);
	nand 	XG12540 	(I23600,g4322,g22360);
	not 	XG12541 	(g20558,I20650);
	and 	XG12542 	(g25125,g23520,g20187);
	and 	XG12543 	(g24725,g23012,g19587);
	and 	XG12544 	(g25112,g23510,g10428);
	or 	XG12545 	(g26703,g10705,g24447);
	or 	XG12546 	(g26770,g10732,g24471);
	or 	XG12547 	(g26737,g10720,g24460);
	and 	XG12548 	(g25371,I24524,g22173,g5062);
	and 	XG12549 	(g24642,g22898,g8290);
	not 	XG12550 	(g21177,I20957);
	and 	XG12551 	(g27281,g26615,g9830);
	and 	XG12552 	(g25420,I24555,g22220,g6058);
	not 	XG12553 	(g20900,I20864);
	nand 	XG12554 	(g25531,g2868,g22763);
	not 	XG12555 	(g20655,I20753);
	and 	XG12556 	(g25110,g23509,g10427);
	nand 	XG12557 	(I22793,I22792,g11956);
	not 	XG12558 	(I22177,g21366);
	not 	XG12559 	(I22180,g21366);
	and 	XG12560 	(g25164,g23569,g16883);
	and 	XG12561 	(g25061,g23461,g17586);
	and 	XG12562 	(g25165,g23570,g14062);
	and 	XG12563 	(g24716,g23004,g15935);
	nand 	XG12564 	(g23786,I22946,I22945);
	not 	XG12565 	(g18882,I19674);
	and 	XG12566 	(g25093,g23493,g12831);
	and 	XG12567 	(g24476,g22330,g18879);
	and 	XG12568 	(g24712,g23001,g19592);
	nand 	XG12569 	(I22800,I22799,g11960);
	and 	XG12570 	(g24998,g23408,g17412);
	nand 	XG12571 	(g25537,g2873,g22763);
	and 	XG12572 	(g25217,g23698,g12418);
	not 	XG12573 	(I22886,g18926);
	not 	XG12574 	(I22889,g18926);
	or 	XG12575 	(g26344,g25010,g2927);
	not 	XG12576 	(g25994,g24575);
	and 	XG12577 	(g25485,I24600,g22220,g6098);
	not 	XG12578 	(g19862,I20233);
	and 	XG12579 	(g24602,g22854,g16507);
	and 	XG12580 	(g24622,g22866,g19856);
	and 	XG12581 	(g24672,g22981,g19534);
	and 	XG12582 	(g24663,g22974,g16621);
	and 	XG12583 	(g24708,g22998,g16474);
	and 	XG12584 	(g24846,I24018,g23555,g3361);
	and 	XG12585 	(g27323,g23086,g26268);
	and 	XG12586 	(g24707,g22997,g13295);
	and 	XG12587 	(g24624,g22867,g16524);
	nor 	XG12588 	(g22513,g19699,g1002);
	nor 	XG12589 	(g22488,g1002,g19699);
	and 	XG12590 	(g24679,g22985,g13289);
	nor 	XG12591 	(g26256,g25479,g23873);
	and 	XG12592 	(g25908,g22520,g24782);
	not 	XG12593 	(g24159,I23321);
	not 	XG12594 	(g24155,I23309);
	not 	XG12595 	(g24154,I23306);
	not 	XG12596 	(g24157,I23315);
	not 	XG12597 	(g24152,I23300);
	not 	XG12598 	(g24158,I23318);
	not 	XG12599 	(g24156,I23312);
	not 	XG12600 	(g24153,I23303);
	not 	XG12601 	(g24160,I23324);
	not 	XG12602 	(g24818,g23191);
	not 	XG12603 	(g22698,I22009);
	and 	XG12604 	(g25510,I24619,g22300,g6444);
	and 	XG12605 	(g25012,g23419,g20644);
	and 	XG12606 	(g24727,g23016,g13300);
	and 	XG12607 	(g24637,g22884,g16586);
	and 	XG12608 	(g25126,g23523,g16839);
	nor 	XG12609 	(g26212,g25408,g23837);
	and 	XG12610 	(g25907,g22519,g24799);
	and 	XG12611 	(g24666,g22975,g11753);
	not 	XG12612 	(g20764,I20819);
	nand 	XG12613 	(I22684,I22683,g11893);
	and 	XG12614 	(g25127,g23524,g13997);
	and 	XG12615 	(g25033,g23433,g17500);
	and 	XG12616 	(g25106,g23506,g17391);
	or 	XG12617 	(g27283,g25924,g25922);
	nand 	XG12618 	(g25779,g24362,g19694);
	and 	XG12619 	(g25014,g23420,g17474);
	and 	XG12620 	(g25166,g23571,g17506);
	and 	XG12621 	(g25071,g23478,g12804);
	and 	XG12622 	(g25040,g23443,g12738);
	or 	XG12623 	(g26894,g18129,g25979);
	and 	XG12624 	(g24668,g22979,g11754);
	and 	XG12625 	(g24635,g22883,g19874);
	not 	XG12626 	(I22785,g18940);
	not 	XG12627 	(I22788,g18940);
	and 	XG12628 	(g25056,g23456,g12779);
	and 	XG12629 	(g25147,g23542,g20202);
	and 	XG12630 	(g25068,g23477,g17574);
	and 	XG12631 	(g24769,g23058,g19619);
	and 	XG12632 	(g25414,I24549,g22194,g5406);
	and 	XG12633 	(g24654,g22922,g11735);
	and 	XG12634 	(g24849,g22227,g4165);
	or 	XG12635 	(g26899,g18199,g26844);
	and 	XG12636 	(g24755,g23030,g16022);
	and 	XG12637 	(g25076,g23479,g12805);
	nand 	XG12638 	(g22663,I21978,I21977);
	or 	XG12639 	(g26673,g10674,g24433);
	nand 	XG12640 	(I22823,I22822,g11978);
	and 	XG12641 	(g25088,g23491,g17601);
	and 	XG12642 	(g24647,g22907,g19903);
	and 	XG12643 	(g24681,g22988,g16653);
	not 	XG12644 	(I22745,g19458);
	not 	XG12645 	(I22748,g19458);
	not 	XG12646 	(g21293,I21036);
	and 	XG12647 	(g24900,I24067,g23582,g3752);
	and 	XG12648 	(g25163,g23566,g20217);
	and 	XG12649 	(g25087,g23489,g17307);
	nand 	XG12650 	(g23810,I22974,I22973);
	and 	XG12651 	(g24709,g23000,g16690);
	not 	XG12652 	(I22557,g20695);
	not 	XG12653 	(I24787,g24266);
	or 	XG12654 	(g26694,g10704,g24444);
	and 	XG12655 	(g25148,g23545,g16867);
	and 	XG12656 	(g24726,g23015,g15965);
	and 	XG12657 	(g24536,g22635,g19516);
	and 	XG12658 	(g26186,g23031,g24580);
	and 	XG12659 	(g27050,g22338,g25789);
	nor 	XG12660 	(g22514,g1018,g19699);
	nor 	XG12661 	(g22448,g19699,g1018);
	and 	XG12662 	(g25043,g23447,g20733);
	and 	XG12663 	(g24861,I24033,g23582,g3712);
	and 	XG12664 	(g25456,I24579,g22210,g5752);
	nand 	XG12665 	(I22894,I22892,g21228);
	nand 	XG12666 	(I22967,I22965,g21228);
	nand 	XG12667 	(I22901,I22899,g21228);
	and 	XG12668 	(g25150,g23547,g17480);
	nor 	XG12669 	(g22539,g19699,g1030);
	nor 	XG12670 	(g22535,g1030,g19699);
	and 	XG12671 	(g25290,I24482,g22173,g5022);
	and 	XG12672 	(g25107,g23508,g17643);
	not 	XG12673 	(g20902,I20870);
	and 	XG12674 	(g25105,g23505,g13973);
	and 	XG12675 	(g24772,g23061,g16287);
	and 	XG12676 	(g25149,g23546,g14030);
	and 	XG12677 	(g27140,g22593,g25885);
	and 	XG12678 	(g25377,I24530,g22210,g5712);
	not 	XG12679 	(g23032,I22211);
	nand 	XG12680 	(I22900,I22899,g12193);
	and 	XG12681 	(g25031,g23432,g20675);
	and 	XG12682 	(g27120,g22543,g25878);
	and 	XG12683 	(g27098,g22528,g25868);
	and 	XG12684 	(g24644,g22903,g11714);
	and 	XG12685 	(g24914,g23301,g8721);
	and 	XG12686 	(g24835,g23233,g8720);
	and 	XG12687 	(g25192,g23648,g20276);
	and 	XG12688 	(g24855,I24027,g23534,g3050);
	and 	XG12689 	(g25086,g23488,g13941);
	and 	XG12690 	(g24822,I24003,g23534,g3010);
	nand 	XG12691 	(g22681,I21994,I21993);
	and 	XG12692 	(g24656,g22926,g11736);
	and 	XG12693 	(g25132,g23528,g10497);
	nand 	XG12694 	(I22966,I22965,g12288);
	and 	XG12695 	(g24754,g23027,g19604);
	nand 	XG12696 	(I22893,I22892,g12189);
	and 	XG12697 	(g25151,g23549,g17719);
	and 	XG12698 	(g24680,g22986,g16422);
	and 	XG12699 	(g24728,g23017,g16513);
	and 	XG12700 	(g25054,g23452,g12778);
	not 	XG12701 	(g21282,I21019);
	and 	XG12702 	(g25178,g23608,g20241);
	not 	XG12703 	(g21246,I20985);
	or 	XG12704 	(g25624,g18224,g24408);
	not 	XG12705 	(I24784,g24265);
	not 	XG12706 	(g21271,I21002);
	nand 	XG12707 	(I23585,g4332,g22409);
	or 	XG12708 	(g27290,g25928,g25926);
	and 	XG12709 	(g25129,g23527,g17682);
	and 	XG12710 	(g25128,g23525,g17418);
	not 	XG12711 	(I22989,g21175);
	nand 	XG12712 	(I23969,g490,g22202);
	and 	XG12713 	(g24684,g22989,g11769);
	and 	XG12714 	(g25079,g23483,g21011);
	not 	XG12715 	(I25356,g24374);
	and 	XG12716 	(g24812,g22192,g19662);
	and 	XG12717 	(g28570,g20434,g27456);
	and 	XG12718 	(g26130,g19772,g24890);
	and 	XG12719 	(g24558,g19566,g22516);
	and 	XG12720 	(g24552,g19538,g22487);
	and 	XG12721 	(g27230,g19558,g25906);
	and 	XG12722 	(g25931,g19477,g24574);
	nand 	XG12723 	(I22711,I22710,g11915);
	or 	XG12724 	(g25622,g18217,g24546);
	and 	XG12725 	(g27300,g26672,g12370);
	and 	XG12726 	(g27292,g26654,g1714);
	or 	XG12727 	(g27563,g24704,g26104);
	and 	XG12728 	(g27340,g26784,g10199);
	or 	XG12729 	(g25633,g18282,g24420);
	nor 	XG12730 	(g22357,g19699,g1024);
	nor 	XG12731 	(g22522,g1024,g19699);
	or 	XG12732 	(g23162,I22267,g20170,g20184);
	and 	XG12733 	(g27293,g26655,g9972);
	or 	XG12734 	(g28089,g18731,g27269);
	or 	XG12735 	(g25894,g23229,g24817);
	or 	XG12736 	(g26912,g18209,g25946);
	and 	XG12737 	(g25921,g9664,g24936);
	and 	XG12738 	(g26094,g9664,g24936);
	and 	XG12739 	(g25915,g9602,g24926);
	and 	XG12740 	(g26084,g9602,g24926);
	or 	XG12741 	(g26898,g18194,g26387);
	or 	XG12742 	(g28088,g18729,g27264);
	nor 	XG12743 	(g22521,g19699,g1036);
	and 	XG12744 	(g25067,g22885,g4722);
	or 	XG12745 	(g23721,I22852,g21385,g21401);
	and 	XG12746 	(g25084,g22885,g4737);
	or 	XG12747 	(g27596,g24775,g26207);
	or 	XG12748 	(g28086,g18702,g27268);
	or 	XG12749 	(g26334,g24591,g1171);
	or 	XG12750 	(g26342,g24591,g8407);
	nand 	XG12751 	(g24880,g22839,g23266,g23281);
	or 	XG12752 	(g28090,g18733,g27275);
	and 	XG12753 	(g25103,g22908,g4927);
	and 	XG12754 	(g27333,g26765,g10180);
	nand 	XG12755 	(g24584,g22715,g22836,g22852);
	nand 	XG12756 	(g24547,g22754,g22643,g22638);
	or 	XG12757 	(g28084,g18698,g27254);
	and 	XG12758 	(g27329,g26743,g12052);
	or 	XG12759 	(g27590,g24764,g26179);
	and 	XG12760 	(g25124,g22908,g4917);
	nor 	XG12761 	(g25950,g24591,g1070);
	nor 	XG12762 	(g25954,g24591,g7750);
	or 	XG12763 	(g23751,I22880,g21402,g21415);
	and 	XG12764 	(g27633,g25766,g13076);
	nor 	XG12765 	(g22545,g19720,g1373);
	nor 	XG12766 	(g22540,g1373,g19720);
	and 	XG12767 	(g26822,g13116,g24841);
	nand 	XG12768 	(g19854,I20223,I20222);
	not 	XG12769 	(g22332,I21838);
	nand 	XG12770 	(g24566,g22713,g22755);
	or 	XG12771 	(g23184,I22280,g20185,g20198);
	or 	XG12772 	(g24254,g18306,g23265);
	nand 	XG12773 	(I22938,I22936,g21228);
	nand 	XG12774 	(I22846,I22844,g21228);
	nand 	XG12775 	(I22873,I22871,g21228);
	nand 	XG12776 	(I22866,I22864,g21228);
	nand 	XG12777 	(I22931,I22929,g21228);
	nand 	XG12778 	(g19782,I20189,I20188);
	nand 	XG12779 	(g24678,g23010,g22994);
	or 	XG12780 	(g26759,g7511,g24468);
	and 	XG12781 	(g27324,g26720,g10150);
	or 	XG12782 	(g26927,g18539,g26711);
	or 	XG12783 	(g26933,g18551,g26808);
	and 	XG12784 	(g27301,g26679,g11992);
	or 	XG12785 	(g28045,g18141,g27378);
	or 	XG12786 	(g26725,g10719,g24457);
	nand 	XG12787 	(g19764,I20167,I20166);
	or 	XG12788 	(g26934,g18556,g26845);
	not 	XG12789 	(g22957,I22143);
	not 	XG12790 	(g22626,I21941);
	or 	XG12791 	(g26328,g24591,g1183);
	or 	XG12792 	(g26327,g24591,g8462);
	and 	XG12793 	(g27305,g26683,g10041);
	nor 	XG12794 	(g22491,g19720,g1361);
	nor 	XG12795 	(g22524,g1361,g19720);
	nand 	XG12796 	(g19792,I20205,I20204);
	nand 	XG12797 	(g24652,g22757,g22940,g22712);
	or 	XG12798 	(g28085,g18700,g27263);
	nand 	XG12799 	(I22754,I22753,g11937);
	not 	XG12800 	(g25423,I24558);
	or 	XG12801 	(g24238,g18248,g23254);
	and 	XG12802 	(g27326,g26731,g12048);
	and 	XG12803 	(g25123,g22885,g4732);
	and 	XG12804 	(g25143,g22908,g4922);
	and 	XG12805 	(g26712,g24463,g24508);
	and 	XG12806 	(g26749,g23578,g24494);
	and 	XG12807 	(g26750,g24474,g24514);
	and 	XG12808 	(g26779,g23620,g24497);
	or 	XG12809 	(g28083,g18689,g27249);
	nand 	XG12810 	(g24544,g22651,g22661,g22666);
	nand 	XG12811 	(g24661,g22984,g23195,g23210);
	or 	XG12812 	(g26931,g18547,g26778);
	or 	XG12813 	(g26932,g18549,g26684);
	and 	XG12814 	(g25085,g22908,g4912);
	or 	XG12815 	(g28087,g18720,g27255);
	not 	XG12816 	(g22976,I22149);
	or 	XG12817 	(g27561,g24702,g26100);
	or 	XG12818 	(g26930,g18544,g26799);
	and 	XG12819 	(g27314,g26702,g12436);
	and 	XG12820 	(g27304,g26682,g2273);
	not 	XG12821 	(g26081,g24619);
	not 	XG12822 	(g25882,g25026);
	not 	XG12823 	(g25899,g24997);
	and 	XG12824 	(g25159,g22908,g4907);
	or 	XG12825 	(g28369,g25938,g27160);
	and 	XG12826 	(g27350,g26803,g10217);
	or 	XG12827 	(g25614,g18161,g24797);
	or 	XG12828 	(g27289,g25927,g25925);
	nor 	XG12829 	(g25947,g24591,g1199);
	nor 	XG12830 	(g25944,g24591,g7716);
	or 	XG12831 	(g27562,g24703,g26102);
	or 	XG12832 	(g26897,g18176,g26611);
	or 	XG12833 	(g26919,g18267,g25951);
	or 	XG12834 	(g26929,g18543,g26635);
	or 	XG12835 	(g26928,g18541,g26713);
	nand 	XG12836 	(I22865,I22864,g12146);
	or 	XG12837 	(g25631,g18275,g24554);
	or 	XG12838 	(g26896,g18171,g26341);
	nand 	XG12839 	(I22718,I22717,g11916);
	or 	XG12840 	(g26793,g7520,g24478);
	or 	XG12841 	(g27551,g24675,g26091);
	or 	XG12842 	(g27589,g24763,g26177);
	or 	XG12843 	(g27579,g24748,g26157);
	and 	XG12844 	(g25102,g22885,g4727);
	or 	XG12845 	(g27569,g24721,g26124);
	nand 	XG12846 	(I22762,I22760,g21434);
	and 	XG12847 	(g25142,g22885,g4717);
	not 	XG12848 	(I26296,g26820);
	nand 	XG12849 	(I22930,I22929,g12223);
	not 	XG12850 	(g23244,I22343);
	not 	XG12851 	(g22546,I21918);
	not 	XG12852 	(g23252,I22353);
	not 	XG12853 	(g23230,I22327);
	not 	XG12854 	(g23219,I22316);
	not 	XG12855 	(g22541,I21911);
	not 	XG12856 	(g23202,I22302);
	not 	XG12857 	(g22592,I21930);
	not 	XG12858 	(g24385,g22908);
	not 	XG12859 	(g24389,g22908);
	not 	XG12860 	(g24404,g22908);
	not 	XG12861 	(g24397,g22908);
	not 	XG12862 	(g24373,g22908);
	not 	XG12863 	(g24384,g22885);
	not 	XG12864 	(g24388,g22885);
	not 	XG12865 	(g24361,g22885);
	not 	XG12866 	(g24396,g22885);
	not 	XG12867 	(g24372,g22885);
	not 	XG12868 	(g25210,g23802);
	not 	XG12869 	(g25244,g23802);
	not 	XG12870 	(g25225,g23802);
	not 	XG12871 	(g25080,g23742);
	not 	XG12872 	(g25197,g23958);
	not 	XG12873 	(g24648,g23148);
	not 	XG12874 	(g25213,g23293);
	not 	XG12875 	(g25032,g23639);
	not 	XG12876 	(g24623,g23076);
	not 	XG12877 	(g25230,g23314);
	not 	XG12878 	(g24527,g22670);
	not 	XG12879 	(g24534,g22670);
	not 	XG12880 	(g24525,g22670);
	not 	XG12881 	(g24516,g22670);
	not 	XG12882 	(g24526,g22942);
	not 	XG12883 	(g24540,g22942);
	not 	XG12884 	(g24535,g22942);
	not 	XG12885 	(g24560,g22942);
	not 	XG12886 	(g24571,g22942);
	not 	XG12887 	(g24548,g22942);
	not 	XG12888 	(g24568,g22942);
	not 	XG12889 	(g24524,g22876);
	not 	XG12890 	(g24533,g22876);
	not 	XG12891 	(g24515,g22689);
	not 	XG12892 	(g24505,g22689);
	not 	XG12893 	(g24509,g22689);
	not 	XG12894 	(g24522,g22689);
	not 	XG12895 	(g24636,g23121);
	not 	XG12896 	(g25264,g23828);
	not 	XG12897 	(g25246,g23828);
	not 	XG12898 	(g25228,g23828);
	not 	XG12899 	(g25044,g23675);
	not 	XG12900 	(g25013,g23599);
	not 	XG12901 	(g25060,g23708);
	and 	XG12902 	(g28238,g19658,g27133);
	and 	XG12903 	(g27351,g26804,g10218);
	nand 	XG12904 	(g27377,g25930,g10685);
	or 	XG12905 	(g26080,g24502,g19393);
	or 	XG12906 	(g26805,g24478,g10776);
	and 	XG12907 	(g28113,g27242,g8016);
	not 	XG12908 	(g28307,g27306);
	and 	XG12909 	(g27363,g26812,g10231);
	and 	XG12910 	(g27723,g21049,g26512);
	and 	XG12911 	(g28304,g19753,g27226);
	nand 	XG12912 	(I22845,I22844,g12113);
	and 	XG12913 	(g27208,g26598,g9037);
	nand 	XG12914 	(g27654,g23042,g26598,g164);
	and 	XG12915 	(g28315,g19769,g27232);
	and 	XG12916 	(g28612,g20539,g27524);
	and 	XG12917 	(g27276,g26607,g9750);
	and 	XG12918 	(g28352,g27705,g10014);
	or 	XG12919 	(g27394,g24573,g25957);
	and 	XG12920 	(g27331,g26754,g10177);
	and 	XG12921 	(g28311,g27679,g9792);
	and 	XG12922 	(g28192,g27415,g8891);
	nand 	XG12923 	(I22761,I22760,g11939);
	and 	XG12924 	(g28630,g20575,g27544);
	and 	XG12925 	(g28554,g20372,g27426);
	and 	XG12926 	(g28587,g20498,g27487);
	nor 	XG12927 	(g25948,g24609,g7752);
	nor 	XG12928 	(g25952,g24609,g1542);
	and 	XG12929 	(g27313,g26701,g1982);
	and 	XG12930 	(g27325,g26724,g12478);
	and 	XG12931 	(g27667,g20601,g26361);
	and 	XG12932 	(g25939,g19490,g24583);
	and 	XG12933 	(g28235,g27592,g9467);
	not 	XG12934 	(g28669,g27705);
	and 	XG12935 	(g27256,g19698,g25937);
	and 	XG12936 	(g25848,g18977,g25539);
	and 	XG12937 	(g27303,g26681,g11996);
	and 	XG12938 	(g27684,g20657,g26386);
	and 	XG12939 	(g27692,g20697,g26392);
	and 	XG12940 	(g28541,g20274,g27403);
	and 	XG12941 	(g28642,g20598,g27555);
	and 	XG12942 	(g27302,g26680,g1848);
	and 	XG12943 	(g27311,g26693,g12431);
	not 	XG12944 	(g27492,g26598);
	and 	XG12945 	(g27676,g20627,g26377);
	and 	XG12946 	(g27316,g26710,g2407);
	and 	XG12947 	(g27328,g26736,g12482);
	and 	XG12948 	(g28555,g20373,g27429);
	and 	XG12949 	(g28569,g20433,g27453);
	and 	XG12950 	(g27315,g26709,g12022);
	and 	XG12951 	(g28601,g20514,g27506);
	nand 	XG12952 	(I22921,g21284,g14677);
	and 	XG12953 	(g27280,g26614,g9825);
	or 	XG12954 	(g27578,g24747,g26155);
	or 	XG12955 	(g27581,g24750,g26161);
	and 	XG12956 	(g28257,g19686,g27179);
	and 	XG12957 	(g27336,g26777,g2675);
	and 	XG12958 	(g27342,g26792,g12592);
	and 	XG12959 	(g27235,g19579,g25910);
	and 	XG12960 	(g28666,g20625,g27567);
	or 	XG12961 	(g27591,g24765,g26181);
	nand 	XG12962 	(I22872,I22871,g12150);
	or 	XG12963 	(g27257,g24498,g25904);
	or 	XG12964 	(g27240,g24467,g25883);
	and 	XG12965 	(g27677,g25888,g13021);
	nor 	XG12966 	(g27046,g25888,g7544);
	nor 	XG12967 	(g25887,g11706,g24984);
	or 	XG12968 	(g27572,g24724,g26129);
	not 	XG12969 	(g27279,g26330);
	nand 	XG12970 	(I22937,I22936,g12226);
	not 	XG12971 	(I25530,g25222);
	and 	XG12972 	(g28330,g19786,g27238);
	or 	XG12973 	(g27570,g24722,g26126);
	and 	XG12974 	(g27284,g26631,g9908);
	and 	XG12975 	(g27330,g26744,g2541);
	and 	XG12976 	(g27334,g26769,g12539);
	and 	XG12977 	(g27312,g26700,g12019);
	and 	XG12978 	(g28258,g19687,g27182);
	and 	XG12979 	(g28706,g20681,g27584);
	and 	XG12980 	(g27560,g20191,g26299);
	and 	XG12981 	(g28247,g19675,g27147);
	and 	XG12982 	(g28602,g20515,g27509);
	and 	XG12983 	(g28333,g19787,g27239);
	and 	XG12984 	(g28248,g19676,g27150);
	and 	XG12985 	(g27699,g20766,g26396);
	not 	XG12986 	(g28620,g27679);
	and 	XG12987 	(g27285,g26632,g9912);
	and 	XG12988 	(g28645,g20599,g27556);
	and 	XG12989 	(g26826,g15747,g24907);
	and 	XG12990 	(g25870,g16182,g24840);
	and 	XG12991 	(g25901,g16290,g24853);
	and 	XG12992 	(g26821,g13103,g24821);
	and 	XG12993 	(g27710,g20904,g26422);
	and 	XG12994 	(g27341,g26788,g10203);
	and 	XG12995 	(g28919,g21295,g27663);
	or 	XG12996 	(g23687,I22830,g21363,g21384);
	and 	XG12997 	(g28627,g20574,g27543);
	and 	XG12998 	(g27616,g20449,g26349);
	and 	XG12999 	(g26633,g20616,g24964);
	and 	XG13000 	(g28346,g19800,g27243);
	not 	XG13001 	(g27018,I25750);
	not 	XG13002 	(I26638,g27965);
	and 	XG13003 	(g28689,g20651,g27575);
	or 	XG13004 	(g27974,g25063,g26544);
	or 	XG13005 	(g27580,g24749,g26159);
	and 	XG13006 	(g27335,g26776,g12087);
	and 	XG13007 	(g28686,g20650,g27574);
	nand 	XG13008 	(g24620,g22874,g22902);
	and 	XG13009 	(g28663,g20624,g27566);
	and 	XG13010 	(g28318,g19770,g27233);
	or 	XG13011 	(g27970,g25050,g26514);
	not 	XG13012 	(g27014,g25888);
	and 	XG13013 	(g28269,g19712,g27205);
	and 	XG13014 	(g28586,g20497,g27484);
	and 	XG13015 	(g25865,g18991,g25545);
	not 	XG13016 	(g27349,g26352);
	and 	XG13017 	(g28617,g20552,g27533);
	or 	XG13018 	(g23771,I22912,g21416,g21432);
	or 	XG13019 	(g24279,g15105,g23218);
	and 	XG13020 	(g28299,g27670,g9716);
	nor 	XG13021 	(g27528,g11083,g26352,g8770);
	and 	XG13022 	(g27099,g26352,g14094);
	and 	XG13023 	(g27158,g16645,g26609);
	and 	XG13024 	(g27184,g13756,g26628);
	and 	XG13025 	(g28227,g27583,g9397);
	not 	XG13026 	(g28648,g27693);
	nand 	XG13027 	(g28500,g12323,g27629,g590);
	and 	XG13028 	(g28193,g27629,g8851);
	and 	XG13029 	(g27087,g26284,g13872);
	and 	XG13030 	(g28108,g27237,g7975);
	not 	XG13031 	(g28294,g27295);
	and 	XG13032 	(g28813,g27038,g4104);
	nand 	XG13033 	(g23975,I23120,I23119);
	or 	XG13034 	(g23198,I22298,g20199,g20214);
	and 	XG13035 	(g25873,g16197,g24854);
	and 	XG13036 	(g25905,g16311,g24879);
	and 	XG13037 	(g26828,g15756,g24919);
	or 	XG13038 	(g23796,I22958,g21433,g21462);
	not 	XG13039 	(I26925,g27015);
	and 	XG13040 	(g27286,g26634,g6856);
	and 	XG13041 	(g27294,g26656,g9975);
	and 	XG13042 	(g27277,g14191,g26359);
	or 	XG13043 	(g27515,g13431,g26051);
	nor 	XG13044 	(g27059,g25895,g7577);
	and 	XG13045 	(g27685,g25895,g13032);
	and 	XG13046 	(g28210,g27554,g9229);
	not 	XG13047 	(g28608,g27670);
	or 	XG13048 	(g28118,g26815,g27821);
	nor 	XG13049 	(g25956,g24609,g1413);
	nor 	XG13050 	(g25958,g24609,g7779);
	and 	XG13051 	(g28215,g27565,g9264);
	and 	XG13052 	(g28144,g27020,g4608);
	and 	XG13053 	(g28154,g27306,g8492);
	or 	XG13054 	(g26335,g24609,g1526);
	or 	XG13055 	(g26329,g24609,g8526);
	not 	XG13056 	(g29172,g27020);
	nand 	XG13057 	(g27463,g23204,g26330,g287);
	and 	XG13058 	(g27041,g26330,g8519);
	not 	XG13059 	(g27017,g25895);
	or 	XG13060 	(g27552,g24676,g26092);
	and 	XG13061 	(g27291,g26653,g11969);
	or 	XG13062 	(g26343,g24609,g1514);
	or 	XG13063 	(g26348,g24609,g8466);
	not 	XG13064 	(g28441,g27629);
	or 	XG13065 	(g26099,g22538,g24506);
	and 	XG13066 	(g28159,g27317,g8553);
	and 	XG13067 	(g28324,g27687,g9875);
	and 	XG13068 	(g28339,g27693,g9946);
	and 	XG13069 	(g27646,g25773,g13094);
	nor 	XG13070 	(g27717,g26745,g9492);
	and 	XG13071 	(g27247,g26745,g2759);
	and 	XG13072 	(g28151,g27295,g8426);
	and 	XG13073 	(g28812,g13037,g26972);
	not 	XG13074 	(g27597,g26745);
	and 	XG13075 	(g28117,g27245,g8075);
	not 	XG13076 	(g28321,g27317);
	and 	XG13077 	(g28219,g27573,g9316);
	not 	XG13078 	(g28633,g27687);
	and 	XG13079 	(g24314,g22228,g4515);
	and 	XG13080 	(g24300,g22228,g15123);
	nor 	XG13081 	(g25141,g10334,g22228);
	and 	XG13082 	(g24291,g22550,g18660);
	and 	XG13083 	(g24326,g22228,g4552);
	and 	XG13084 	(g24327,g22228,g4549);
	and 	XG13085 	(g24191,g22722,g319);
	and 	XG13086 	(g24299,g22550,g4456);
	and 	XG13087 	(g24333,g22228,g4512);
	and 	XG13088 	(g24288,g22550,g4417);
	and 	XG13089 	(g24189,g22722,g324);
	nor 	XG13090 	(g25504,g7222,g22550);
	and 	XG13091 	(g24289,g22550,g4427);
	and 	XG13092 	(g24306,g22228,g4483);
	or 	XG13093 	(I25612,g25570,g25569,g25568,g25567);
	or 	XG13094 	(I25613,g25574,g25573,g25572,g25571);
	and 	XG13095 	(g24226,g22594,g446);
	not 	XG13096 	(I25359,g24715);
	and 	XG13097 	(g24190,g22722,g329);
	and 	XG13098 	(g24287,g22550,g4401);
	nand 	XG13099 	(I25219,g24718,g482);
	not 	XG13100 	(g25640,I24781);
	and 	XG13101 	(g24194,g22722,g106);
	and 	XG13102 	(g24324,g22228,g4540);
	and 	XG13103 	(g24301,g22228,g6961);
	and 	XG13104 	(g24197,g22722,g347);
	and 	XG13105 	(g24218,g22594,g872);
	and 	XG13106 	(g24286,g22550,g4405);
	and 	XG13107 	(g24298,g22550,g4392);
	and 	XG13108 	(g24329,g22228,g4462);
	and 	XG13109 	(g24293,g22550,g4438);
	and 	XG13110 	(g24186,g22722,g18102);
	and 	XG13111 	(g24308,g22228,g4489);
	and 	XG13112 	(g24230,g22594,g901);
	and 	XG13113 	(g24323,g22228,g4546);
	and 	XG13114 	(g24316,g22228,g4527);
	and 	XG13115 	(g24319,g22228,g4561);
	and 	XG13116 	(g24229,g22594,g896);
	or 	XG13117 	(g24561,I23756,I23755);
	and 	XG13118 	(g24220,g22594,g255);
	and 	XG13119 	(g24187,g22722,g305);
	and 	XG13120 	(g24193,g22722,g336);
	and 	XG13121 	(g24188,g22722,g316);
	and 	XG13122 	(g24312,g22228,g4501);
	and 	XG13123 	(g24227,g22594,g890);
	and 	XG13124 	(g24302,g22228,g15124);
	and 	XG13125 	(g24295,g22550,g4434);
	and 	XG13126 	(g24292,g22550,g4443);
	and 	XG13127 	(g24228,g22594,g862);
	and 	XG13128 	(g24322,g22228,g4423);
	and 	XG13129 	(g24195,g22722,g74);
	and 	XG13130 	(g24330,g22228,g18661);
	and 	XG13131 	(g24222,g22594,g262);
	and 	XG13132 	(g24309,g22228,g4480);
	and 	XG13133 	(g24304,g22228,g12875);
	and 	XG13134 	(g24283,g22550,g4411);
	and 	XG13135 	(g24224,g22594,g269);
	and 	XG13136 	(g24196,g22722,g333);
	and 	XG13137 	(g24297,g22550,g4455);
	and 	XG13138 	(g24221,g22594,g232);
	and 	XG13139 	(g24320,g22228,g6973);
	and 	XG13140 	(g24290,g22550,g4430);
	and 	XG13141 	(g24285,g22550,g4388);
	and 	XG13142 	(g24332,g22228,g4459);
	or 	XG13143 	(g25694,g18738,g24638);
	and 	XG13144 	(g24303,g22228,g4369);
	not 	XG13145 	(I25327,g24641);
	and 	XG13146 	(g24313,g22228,g4504);
	and 	XG13147 	(g24307,g22228,g4486);
	and 	XG13148 	(g24219,g22594,g225);
	and 	XG13149 	(g24294,g22550,g4452);
	and 	XG13150 	(g24223,g22594,g239);
	and 	XG13151 	(g24311,g22228,g4498);
	or 	XG13152 	(g25693,g18707,g24627);
	and 	XG13153 	(g24225,g22594,g246);
	and 	XG13154 	(g24217,g22594,g18200);
	and 	XG13155 	(g24199,g22722,g355);
	and 	XG13156 	(g24310,g22228,g4495);
	and 	XG13157 	(g24296,g22550,g4382);
	and 	XG13158 	(g24198,g22722,g351);
	and 	XG13159 	(g24317,g22228,g4534);
	and 	XG13160 	(g24325,g22228,g4543);
	and 	XG13161 	(g24305,g22228,g4477);
	and 	XG13162 	(g24284,g22550,g4375);
	and 	XG13163 	(g24331,g22228,g6977);
	and 	XG13164 	(g24321,g22228,g4558);
	and 	XG13165 	(g24315,g22228,g4521);
	and 	XG13166 	(g24328,g22228,g4567);
	and 	XG13167 	(g24192,g22722,g311);
	nand 	XG13168 	(I25242,g24744,g490);
	and 	XG13169 	(g24318,g22228,g4555);
	not 	XG13170 	(g24893,I24060);
	not 	XG13171 	(g24866,I24038);
	not 	XG13172 	(g25064,I24228);
	not 	XG13173 	(g24920,I24089);
	not 	XG13174 	(g24911,I24078);
	not 	XG13175 	(g25051,I24215);
	not 	XG13176 	(g25027,I24191);
	not 	XG13177 	(g24869,I24041);
	not 	XG13178 	(g24850,I24022);
	not 	XG13179 	(g24836,I24008);
	not 	XG13180 	(g24819,I23998);
	or 	XG13181 	(g27008,I25736,g21370,g26866);
	nor 	XG13182 	(g27511,g20277,g26866,g22137);
	not 	XG13183 	(g25250,I24434);
	not 	XG13184 	(g24490,g22594);
	not 	XG13185 	(g24366,g22594);
	not 	XG13186 	(g24377,g22594);
	not 	XG13187 	(g24407,g22594);
	not 	XG13188 	(g25563,g22594);
	not 	XG13189 	(g24365,g22594);
	not 	XG13190 	(g25538,g22594);
	not 	XG13191 	(g24386,g22594);
	not 	XG13192 	(g24356,g22594);
	not 	XG13193 	(g25544,g22594);
	not 	XG13194 	(g25558,g22594);
	not 	XG13195 	(g25528,g22594);
	not 	XG13196 	(g25552,g22594);
	not 	XG13197 	(g24426,g22722);
	not 	XG13198 	(g24376,g22722);
	not 	XG13199 	(g24438,g22722);
	not 	XG13200 	(g24418,g22722);
	not 	XG13201 	(g24419,g22722);
	not 	XG13202 	(g24424,g22722);
	not 	XG13203 	(g24364,g22722);
	not 	XG13204 	(g24425,g22722);
	not 	XG13205 	(g24375,g22722);
	not 	XG13206 	(g24428,g22722);
	not 	XG13207 	(g24429,g22722);
	not 	XG13208 	(g24405,g22722);
	not 	XG13209 	(g24452,g22722);
	not 	XG13210 	(g24431,g22722);
	not 	XG13211 	(g25553,g22550);
	not 	XG13212 	(g24367,g22550);
	not 	XG13213 	(g25523,g22550);
	not 	XG13214 	(g24358,g22550);
	not 	XG13215 	(g24359,g22550);
	not 	XG13216 	(g25546,g22550);
	not 	XG13217 	(g25547,g22550);
	not 	XG13218 	(g24379,g22550);
	not 	XG13219 	(g25554,g22550);
	not 	XG13220 	(g25566,g22550);
	not 	XG13221 	(g25555,g22550);
	not 	XG13222 	(g25560,g22550);
	not 	XG13223 	(g25525,g22550);
	not 	XG13224 	(g25561,g22550);
	not 	XG13225 	(g25533,g22550);
	not 	XG13226 	(g25548,g22550);
	not 	XG13227 	(g25452,g22228);
	not 	XG13228 	(g25326,g22228);
	not 	XG13229 	(g25409,g22228);
	not 	XG13230 	(g24394,g22228);
	not 	XG13231 	(g24360,g22228);
	not 	XG13232 	(g25517,g22228);
	not 	XG13233 	(g25410,g22228);
	not 	XG13234 	(g25286,g22228);
	not 	XG13235 	(g25287,g22228);
	not 	XG13236 	(g25480,g22228);
	not 	XG13237 	(g25231,g22228);
	not 	XG13238 	(g25481,g22228);
	not 	XG13239 	(g25370,g22228);
	not 	XG13240 	(g25451,g22228);
	not 	XG13241 	(g25140,g22228);
	not 	XG13242 	(g25324,g22228);
	not 	XG13243 	(g25506,g22228);
	not 	XG13244 	(g25325,g22228);
	not 	XG13245 	(g25214,g22228);
	not 	XG13246 	(g24368,g22228);
	not 	XG13247 	(g25185,g22228);
	not 	XG13248 	(g25524,g22228);
	not 	XG13249 	(g25266,g22228);
	not 	XG13250 	(g25267,g22228);
	not 	XG13251 	(g25288,g22228);
	not 	XG13252 	(g25289,g22228);
	not 	XG13253 	(g25158,g22228);
	not 	XG13254 	(g25171,g22228);
	not 	XG13255 	(g25198,g22228);
	not 	XG13256 	(g25232,g22228);
	not 	XG13257 	(g25369,g22228);
	not 	XG13258 	(g25505,g22228);
	not 	XG13259 	(g25248,g22228);
	not 	XG13260 	(g25249,g22228);
	and 	XG13261 	(g28677,g20635,g27571);
	and 	XG13262 	(g28451,g20090,g27283);
	and 	XG13263 	(g28456,g20104,g27290);
	or 	XG13264 	(g25688,g21887,g24812);
	not 	XG13265 	(g26424,I25356);
	nand 	XG13266 	(I23986,I23985,g22182);
	nand 	XG13267 	(I23601,I23600,g22360);
	nand 	XG13268 	(I23586,I23585,g22409);
	nand 	XG13269 	(I23970,I23969,g22202);
	or 	XG13270 	(g25752,g22099,g25079);
	or 	XG13271 	(g25677,g21834,g24684);
	nand 	XG13272 	(g23575,I22712,I22711);
	nand 	XG13273 	(g24933,g23154,g19466);
	nand 	XG13274 	(g24972,g23172,g19962);
	nand 	XG13275 	(I23971,I23969,g490);
	nand 	XG13276 	(g24943,g23172,g20068);
	not 	XG13277 	(g23823,I22989);
	nand 	XG13278 	(g25019,g23172,g20055);
	or 	XG13279 	(g25731,g22014,g25128);
	or 	XG13280 	(g25744,g22059,g25129);
	nand 	XG13281 	(g24958,g23462,g21330);
	nand 	XG13282 	(g25021,g23363,g21417);
	or 	XG13283 	(g28077,g21879,g27120);
	nand 	XG13284 	(I23587,I23585,g4332);
	or 	XG13285 	(g26940,g21886,g25908);
	or 	XG13286 	(g25742,g22057,g25093);
	nand 	XG13287 	(g24989,g23363,g21345);
	not 	XG13288 	(g23824,g21271);
	not 	XG13289 	(g25641,I24784);
	or 	XG13290 	(g28043,g21714,g27323);
	not 	XG13291 	(g23800,g21246);
	or 	XG13292 	(g25741,g22056,g25178);
	not 	XG13293 	(I22576,g21282);
	or 	XG13294 	(g25701,g21920,g25054);
	nand 	XG13295 	(g25002,g23154,g19474);
	or 	XG13296 	(g27858,g26737,g17405);
	or 	XG13297 	(g27800,g26703,g17321);
	or 	XG13298 	(g25679,g21836,g24728);
	nand 	XG13299 	(g24942,g23172,g20039);
	nand 	XG13300 	(g24934,g23462,g21283);
	or 	XG13301 	(g25650,g21743,g24663);
	or 	XG13302 	(g25651,g21744,g24680);
	or 	XG13303 	(g25759,g22106,g25166);
	or 	XG13304 	(g25758,g22105,g25151);
	nand 	XG13305 	(g23761,I22894,I22893);
	nand 	XG13306 	(g24917,g23172,g19913);
	or 	XG13307 	(g25661,g21786,g24754);
	nand 	XG13308 	(g23809,I22967,I22966);
	or 	XG13309 	(g25757,g22104,g25132);
	or 	XG13310 	(g25662,g21787,g24656);
	or 	XG13311 	(g26939,g21884,g25907);
	and 	XG13312 	(g24688,g22663,g22681);
	nor 	XG13313 	(g26515,g24822,g24843);
	or 	XG13314 	(g26616,g24822,g24843,g24855,g24881);
	or 	XG13315 	(g25730,g22013,g25107);
	or 	XG13316 	(g28078,g21880,g27140);
	or 	XG13317 	(g25698,g21917,g25104);
	or 	XG13318 	(g25697,g21916,g25086);
	or 	XG13319 	(g25592,g21706,g24672);
	or 	XG13320 	(g25649,g21742,g24654);
	nor 	XG13321 	(g26545,g24855,g24881);
	or 	XG13322 	(g28578,g26273,g27327);
	or 	XG13323 	(g25755,g22102,g25192);
	or 	XG13324 	(g25595,g21717,g24835);
	or 	XG13325 	(g25599,g21721,g24914);
	or 	XG13326 	(g25648,g21741,g24644);
	or 	XG13327 	(g28076,g21878,g27098);
	or 	XG13328 	(g28075,g21877,g27083);
	or 	XG13329 	(g25710,g21961,g25031);
	or 	XG13330 	(g25695,g21914,g24998);
	nand 	XG13331 	(g23762,I22901,I22900);
	or 	XG13332 	(g25678,g21835,g24709);
	or 	XG13333 	(g28518,g26158,g27281);
	nand 	XG13334 	(g24924,g23172,g20007);
	nor 	XG13335 	(g25770,g25377,g25417);
	or 	XG13336 	(g25821,g25377,g25417,g25456,g25482);
	nand 	XG13337 	(g25532,g23363,g21360);
	or 	XG13338 	(g25739,g22054,g25149);
	or 	XG13339 	(g25740,g22055,g25164);
	or 	XG13340 	(g25594,g21708,g24772);
	or 	XG13341 	(g25712,g21963,g25126);
	or 	XG13342 	(g25711,g21962,g25105);
	not 	XG13343 	(g23746,g20902);
	nor 	XG13344 	(g26865,g25290,g25328);
	or 	XG13345 	(g25791,g25290,g25328,g25371,g25411);
	or 	XG13346 	(g27907,g26770,g17424);
	or 	XG13347 	(g25745,g22060,g25150);
	nor 	XG13348 	(g25777,g25456,g25482);
	or 	XG13349 	(g25729,g22012,g25091);
	nor 	XG13350 	(g26574,g24861,g24887);
	or 	XG13351 	(g26657,g24861,g24887,g24900,g24908);
	and 	XG13352 	(g25223,g10652,g22523);
	or 	XG13353 	(g24518,g7601,g22517);
	or 	XG13354 	(g25724,g22007,g25043);
	or 	XG13355 	(g25728,g22011,g25076);
	or 	XG13356 	(g25690,g21889,g24864);
	or 	XG13357 	(g28070,g21867,g27050);
	or 	XG13358 	(g26938,g21883,g26186);
	or 	XG13359 	(g25691,g21890,g24536);
	or 	XG13360 	(g25660,g21785,g24726);
	or 	XG13361 	(g25726,g22009,g25148);
	or 	XG13362 	(g25727,g22010,g25163);
	and 	XG13363 	(g27265,g26759,g26785);
	and 	XG13364 	(g27614,g26759,g26785);
	and 	XG13365 	(g27251,g26694,g26721);
	and 	XG13366 	(g27594,g26694,g26721);
	not 	XG13367 	(g27975,g26694);
	not 	XG13368 	(g27088,g26694);
	not 	XG13369 	(g25642,I24787);
	not 	XG13370 	(g23440,I22557);
	or 	XG13371 	(g25700,g21919,g25040);
	and 	XG13372 	(g25357,g23786,g23810);
	or 	XG13373 	(g25702,g21921,g25068);
	or 	XG13374 	(g25703,g21922,g25087);
	nor 	XG13375 	(g26603,g24900,g24908);
	nand 	XG13376 	(g24918,g23088,g136);
	not 	XG13377 	(g23870,g21293);
	not 	XG13378 	(g23613,I22748);
	or 	XG13379 	(g25665,g21790,g24708);
	or 	XG13380 	(g25664,g21789,g24681);
	or 	XG13381 	(g25672,g21829,g24647);
	or 	XG13382 	(g25716,g21967,g25088);
	nand 	XG13383 	(g23685,I22824,I22823);
	nand 	XG13384 	(g25003,g23462,g21353);
	and 	XG13385 	(g27600,g26725,g26755);
	and 	XG13386 	(g27259,g26725,g26755);
	and 	XG13387 	(g27246,g26673,g26690);
	and 	XG13388 	(g27588,g26673,g26690);
	not 	XG13389 	(g27971,g26673);
	not 	XG13390 	(g27084,g26673);
	and 	XG13391 	(g25207,g10621,g22513);
	or 	XG13392 	(g24510,g7567,g22488);
	or 	XG13393 	(g25666,g21793,g24788);
	or 	XG13394 	(g25676,g21833,g24668);
	or 	XG13395 	(g25674,g21831,g24755);
	or 	XG13396 	(g25675,g21832,g24769);
	or 	XG13397 	(g25689,g21888,g24849);
	nor 	XG13398 	(g25769,g25414,g25453);
	or 	XG13399 	(g25805,g25331,g25374,g25414,g25453);
	or 	XG13400 	(g25715,g21966,g25071);
	or 	XG13401 	(g25713,g21964,g25147);
	nand 	XG13402 	(g24957,g23462,g21359);
	or 	XG13403 	(g25717,g21968,g25106);
	or 	XG13404 	(g25723,g22006,g25033);
	or 	XG13405 	(g25714,g21965,g25056);
	not 	XG13406 	(g23653,I22788);
	or 	XG13407 	(g25658,g21783,g24635);
	nand 	XG13408 	(g25381,g23088,g538);
	or 	XG13409 	(g25737,g22052,g25045);
	nand 	XG13410 	(g25048,g23088,g542);
	or 	XG13411 	(g25709,g21960,g25014);
	nand 	XG13412 	(g23616,I22755,I22754);
	or 	XG13413 	(g25671,g21828,g24637);
	or 	XG13414 	(g25725,g22008,g25127);
	nand 	XG13415 	(g23552,I22685,I22684);
	not 	XG13416 	(g23715,g20764);
	nand 	XG13417 	(g24916,g23154,g19450);
	or 	XG13418 	(g25663,g21788,g24666);
	nand 	XG13419 	(I25845,g24799,g26212);
	or 	XG13420 	(g25685,g21866,g24476);
	or 	XG13421 	(g28073,g21875,g27097);
	or 	XG13422 	(g25673,g21830,g24727);
	nand 	XG13423 	(g24951,g23088,g199);
	or 	XG13424 	(g25696,g21915,g25012);
	nand 	XG13425 	(g25049,g23462,g21344);
	nor 	XG13426 	(g25800,g25510,g25518);
	or 	XG13427 	(g25856,g25462,g25488,g25510,g25518);
	not 	XG13428 	(g26337,g24818);
	nand 	XG13429 	(g25038,g23363,g21331);
	nand 	XG13430 	(I25907,g24782,g26256);
	nand 	XG13431 	(g24906,g23088,g8743);
	or 	XG13432 	(g25645,g21738,g24679);
	or 	XG13433 	(g25646,g21739,g24706);
	nand 	XG13434 	(g25425,g23172,g20081);
	or 	XG13435 	(g25597,g21719,g24892);
	or 	XG13436 	(g25657,g21782,g24624);
	or 	XG13437 	(g25659,g21784,g24707);
	nor 	XG13438 	(g26546,g24846,g24858);
	or 	XG13439 	(g26636,g24846,g24858,g24884,g24897);
	nand 	XG13440 	(g24974,g23363,g21301);
	or 	XG13441 	(g25746,g22063,g25217);
	or 	XG13442 	(g25644,g21737,g24622);
	or 	XG13443 	(g25643,g21736,g24602);
	not 	XG13444 	(I22816,g19862);
	not 	XG13445 	(I22819,g19862);
	nor 	XG13446 	(g25784,g25485,g25507);
	or 	XG13447 	(g25839,g25420,g25459,g25485,g25507);
	or 	XG13448 	(g25743,g22058,g25110);
	or 	XG13449 	(g25593,g21707,g24716);
	nand 	XG13450 	(g24944,g23363,g21354);
	not 	XG13451 	(g27585,g25994);
	nand 	XG13452 	(g25020,g23462,g21377);
	not 	XG13453 	(g23760,I22889);
	nand 	XG13454 	(g24975,g23363,g21388);
	nand 	XG13455 	(g24932,g23172,g19886);
	or 	XG13456 	(g25756,g22103,g25112);
	not 	XG13457 	(I25586,g25537);
	nand 	XG13458 	(g23656,I22801,I22800);
	or 	XG13459 	(g25686,g21881,g24712);
	nand 	XG13460 	(g24925,g23154,g20092);
	or 	XG13461 	(g25751,g22098,g25061);
	not 	XG13462 	(g22171,g18882);
	nand 	XG13463 	(g25018,g23154,g20107);
	or 	XG13464 	(g25591,g21705,g24642);
	nand 	XG13465 	(g25062,g23363,g21403);
	or 	XG13466 	(g25753,g22100,g25165);
	or 	XG13467 	(g25760,g22109,g25238);
	not 	XG13468 	(g23003,I22180);
	nand 	XG13469 	(g23655,I22794,I22793);
	not 	XG13470 	(g23651,g20655);
	not 	XG13471 	(I25594,g25531);
	not 	XG13472 	(g23745,g20900);
	nand 	XG13473 	(g23576,I22719,I22718);
	nor 	XG13474 	(g25778,g25420,g25459);
	not 	XG13475 	(g23776,g21177);
	or 	XG13476 	(g25754,g22101,g25179);
	nor 	XG13477 	(g26872,g25371,g25411);
	and 	XG13478 	(g27601,g26737,g26766);
	and 	XG13479 	(g27260,g26737,g26766);
	not 	XG13480 	(g27092,g26737);
	not 	XG13481 	(g27984,g26737);
	and 	XG13482 	(g27266,g26770,g26789);
	and 	XG13483 	(g27615,g26770,g26789);
	not 	XG13484 	(g27990,g26770);
	not 	XG13485 	(g27101,g26770);
	and 	XG13486 	(g27595,g26703,g26733);
	and 	XG13487 	(g27252,g26703,g26733);
	not 	XG13488 	(g27089,g26703);
	not 	XG13489 	(g27976,g26703);
	or 	XG13490 	(g25647,g21740,g24725);
	or 	XG13491 	(g25699,g21918,g25125);
	not 	XG13492 	(g23529,g20558);
	nand 	XG13493 	(I23602,I23600,g4322);
	nand 	XG13494 	(g25527,g23462,g21294);
	or 	XG13495 	(g25704,g21925,g25173);
	not 	XG13496 	(I24445,g22923);
	not 	XG13497 	(I24448,g22923);
	or 	XG13498 	(g28071,g21873,g27085);
	or 	XG13499 	(g28072,g21874,g27086);
	or 	XG13500 	(g25738,g22053,g25059);
	or 	XG13501 	(g25596,g21718,g24865);
	or 	XG13502 	(g28074,g21876,g27119);
	nand 	XG13503 	(g24950,g23154,g19442);
	or 	XG13504 	(g28591,g26286,g27332);
	or 	XG13505 	(I24117,g23172,g23154,g23088);
	or 	XG13506 	(g25598,g21720,g24904);
	nor 	XG13507 	(g25785,g25462,g25488);
	nor 	XG13508 	(g26573,g24884,g24897);
	not 	XG13509 	(g23650,g20653);
	or 	XG13510 	(g25687,g21882,g24729);
	or 	XG13511 	(g25732,g22017,g25201);
	or 	XG13512 	(g25718,g21971,g25187);
	or 	XG13513 	(g25652,g21747,g24777);
	and 	XG13514 	(g26484,g8841,g24946);
	and 	XG13515 	(g26398,g10474,g24946);
	or 	XG13516 	(g25680,g21839,g24794);
	nor 	XG13517 	(g26873,g25331,g25374);
	not 	XG13518 	(g23231,g20050);
	and 	XG13519 	(g24485,g22319,g10710);
	and 	XG13520 	(g24537,g10851,g22626);
	and 	XG13521 	(g24541,g10851,g22626);
	and 	XG13522 	(g24491,g22332,g10727);
	and 	XG13523 	(g24872,g9104,g23088);
	or 	XG13524 	(g28544,g26229,g27300);
	nand 	XG13525 	(g24905,g23088,g534);
	and 	XG13526 	(g27634,g26793,g26805);
	and 	XG13527 	(g27270,g26793,g26805);
	not 	XG13528 	(I24497,g22592);
	not 	XG13529 	(I23671,g23202);
	not 	XG13530 	(I24455,g22541);
	not 	XG13531 	(I23680,g23219);
	not 	XG13532 	(I23684,g23230);
	not 	XG13533 	(I23694,g23252);
	not 	XG13534 	(I24474,g22546);
	not 	XG13535 	(I23688,g23244);
	and 	XG13536 	(g26485,g10502,g24968);
	and 	XG13537 	(g26516,g8876,g24968);
	nand 	XG13538 	(I23949,g13603,g23162);
	nand 	XG13539 	(g23719,I22846,I22845);
	nand 	XG13540 	(g24988,g23088,g546);
	nand 	XG13541 	(g23780,I22931,I22930);
	nand 	XG13542 	(g24973,g23462,g21272);
	nand 	XG13543 	(g23617,I22762,I22761);
	or 	XG13544 	(g28534,g26204,g27292);
	not 	XG13545 	(g27662,I26296);
	and 	XG13546 	(g27598,g10475,g25899);
	and 	XG13547 	(g27648,g8974,g25882);
	nand 	XG13548 	(I23987,I23985,g482);
	not 	XG13549 	(g27994,g26793);
	not 	XG13550 	(g27112,g26793);
	nand 	XG13551 	(I24383,g14347,g23721);
	or 	XG13552 	(g25632,g18277,g24558);
	nand 	XG13553 	(g23747,I22866,I22865);
	or 	XG13554 	(g28564,g26252,g27314);
	or 	XG13555 	(g28545,g26230,g27301);
	or 	XG13556 	(g28536,g26205,g27293);
	or 	XG13557 	(g28056,g18210,g27230);
	and 	XG13558 	(g27958,g22449,g25950);
	and 	XG13559 	(g27962,g19597,g25954);
	nand 	XG13560 	(g24567,g2917,g22957);
	nand 	XG13561 	(g23748,I22873,I22872);
	or 	XG13562 	(g28613,g26310,g27350);
	or 	XG13563 	(g28577,g26272,g27326);
	nand 	XG13564 	(g24621,g2927,g22957);
	not 	XG13565 	(g27576,g26081);
	or 	XG13566 	(g28549,g26233,g27304);
	or 	XG13567 	(g26944,g18658,g26130);
	not 	XG13568 	(I24334,g22976);
	not 	XG13569 	(I24331,g22976);
	nand 	XG13570 	(g23781,I22938,I22937);
	nor 	XG13571 	(g27102,g26779,g26750);
	nor 	XG13572 	(g27093,g26749,g26712);
	nand 	XG13573 	(g24601,g2965,g22957);
	or 	XG13574 	(g27019,g14610,g26822);
	and 	XG13575 	(g24929,g20875,g23751);
	and 	XG13576 	(g27025,g7917,g26334);
	and 	XG13577 	(g27028,g1157,g26342);
	or 	XG13578 	(g27742,g26673,g17292);
	not 	XG13579 	(I25190,g25423);
	or 	XG13580 	(g27779,g26694,g17317);
	nor 	XG13581 	(g24631,g22957,g20219,g20436,g20516);
	not 	XG13582 	(g27091,g26725);
	not 	XG13583 	(g27983,g26725);
	nand 	XG13584 	(I24414,g14382,g23751);
	or 	XG13585 	(g29293,g18777,g28570);
	not 	XG13586 	(g27100,g26759);
	not 	XG13587 	(g27989,g26759);
	and 	XG13588 	(g28165,g22455,g27018);
	or 	XG13589 	(g28581,g26276,g27329);
	or 	XG13590 	(g25960,g24678,g24566);
	or 	XG13591 	(g25623,g18219,g24552);
	or 	XG13592 	(g28592,g26288,g27333);
	or 	XG13593 	(g26918,g18243,g25931);
	and 	XG13594 	(g24549,g20887,g23162);
	and 	XG13595 	(g28712,g20708,g27590);
	and 	XG13596 	(g28697,g20669,g27581);
	and 	XG13597 	(g28695,g20666,g27580);
	and 	XG13598 	(g28679,g20638,g27572);
	and 	XG13599 	(g28658,g20611,g27563);
	and 	XG13600 	(g22873,g19683,g19854);
	and 	XG13601 	(g22938,g19739,g19782);
	and 	XG13602 	(g28110,g18886,g27974);
	and 	XG13603 	(g28676,g20632,g27570);
	and 	XG13604 	(g28692,g20661,g27578);
	and 	XG13605 	(g28638,g20583,g27551);
	and 	XG13606 	(g28655,g20603,g27561);
	and 	XG13607 	(g22920,g19719,g19764);
	and 	XG13608 	(g22861,g19670,g19792);
	and 	XG13609 	(g28107,g18874,g27970);
	and 	XG13610 	(g28657,g20606,g27562);
	and 	XG13611 	(g28674,g20629,g27569);
	and 	XG13612 	(g28714,g20711,g27591);
	and 	XG13613 	(g28725,g20779,g27596);
	and 	XG13614 	(g29837,g20144,g28369);
	and 	XG13615 	(g28426,g20006,g27257);
	and 	XG13616 	(g27362,g20036,g26080);
	and 	XG13617 	(g28455,g20103,g27289);
	and 	XG13618 	(g28532,g20265,g27394);
	and 	XG13619 	(g28341,g19790,g27240);
	and 	XG13620 	(g28710,g20703,g27589);
	and 	XG13621 	(g28694,g20664,g27579);
	or 	XG13622 	(g28582,g26277,g27330);
	and 	XG13623 	(g26864,g24548,g2907);
	and 	XG13624 	(g28182,g27349,g8770);
	or 	XG13625 	(g28603,g26300,g27340);
	or 	XG13626 	(g28551,g26234,g27305);
	or 	XG13627 	(g29302,g18798,g28601);
	or 	XG13628 	(g29264,g18618,g28248);
	nand 	XG13629 	(I23961,g13631,g23184);
	and 	XG13630 	(g27959,g19374,g25948);
	and 	XG13631 	(g27963,g16047,g25952);
	and 	XG13632 	(g26079,g25060,g6199);
	or 	XG13633 	(g26920,g18283,g25865);
	and 	XG13634 	(g26829,g24505,g2844);
	and 	XG13635 	(g26048,g25044,g5853);
	and 	XG13636 	(g26019,g25032,g5507);
	nand 	XG13637 	(g24662,g2955,g22957);
	or 	XG13638 	(g27278,g25921,g15786);
	or 	XG13639 	(g27542,g26094,g16190);
	or 	XG13640 	(g27532,g26084,g16176);
	or 	XG13641 	(g27274,g25915,g15779);
	and 	XG13642 	(g24921,g20739,g23721);
	or 	XG13643 	(g28052,g18167,g27710);
	and 	XG13644 	(g25866,g24648,g3853);
	or 	XG13645 	(g29282,g18745,g28617);
	or 	XG13646 	(g29283,g18746,g28627);
	nand 	XG13647 	(g28167,g27046,g925);
	and 	XG13648 	(g28558,g27046,g7301);
	nand 	XG13649 	(g24570,g2941,g22957);
	and 	XG13650 	(g24555,g21024,g23184);
	or 	XG13651 	(g29299,g18794,g28587);
	and 	XG13652 	(g25986,g25013,g5160);
	and 	XG13653 	(g25831,g24623,g3151);
	or 	XG13654 	(g26925,g18301,g25939);
	or 	XG13655 	(g29296,g18781,g28586);
	and 	XG13656 	(g27029,g11031,g26327);
	and 	XG13657 	(g27034,g8609,g26328);
	and 	XG13658 	(g26833,g24509,g2852);
	nand 	XG13659 	(g28448,g27377,g23975);
	or 	XG13660 	(g29273,g18639,g28269);
	or 	XG13661 	(g28055,g18190,g27560);
	or 	XG13662 	(g29078,g26572,g27633);
	or 	XG13663 	(g27886,g26759,g14438);
	or 	XG13664 	(g27837,g26725,g17401);
	and 	XG13665 	(g26855,g24535,g2960);
	or 	XG13666 	(g29265,g18620,g28318);
	or 	XG13667 	(g29266,g18621,g28330);
	or 	XG13668 	(g28044,g18130,g27256);
	or 	XG13669 	(g29295,g18780,g28663);
	or 	XG13670 	(g27937,g26793,g14506);
	nand 	XG13671 	(I22922,I22921,g14677);
	nand 	XG13672 	(g24677,g2975,g22957);
	or 	XG13673 	(g29301,g18797,g28686);
	or 	XG13674 	(g29300,g18796,g28666);
	or 	XG13675 	(g28595,g26290,g27335);
	or 	XG13676 	(g29306,g18813,g28689);
	or 	XG13677 	(g29307,g18814,g28706);
	not 	XG13678 	(g28137,I26638);
	or 	XG13679 	(g29272,g18638,g28346);
	and 	XG13680 	(g26301,g25244,g2145);
	or 	XG13681 	(g28574,g26270,g27324);
	or 	XG13682 	(g26926,g18531,g26633);
	or 	XG13683 	(g28060,g18532,g27616);
	or 	XG13684 	(g29284,g18747,g28554);
	or 	XG13685 	(g26913,g18225,g25848);
	and 	XG13686 	(g26088,g25080,g6545);
	or 	XG13687 	(g28580,g26275,g27328);
	or 	XG13688 	(g29224,g18156,g28919);
	and 	XG13689 	(g26274,g25210,g2130);
	or 	XG13690 	(g28576,g26271,g27325);
	nand 	XG13691 	(g24576,g2902,g22957);
	or 	XG13692 	(g29270,g18635,g28258);
	or 	XG13693 	(g28548,g26232,g27303);
	or 	XG13694 	(g28605,g26302,g27341);
	or 	XG13695 	(g28054,g18170,g27723);
	and 	XG13696 	(g28204,g27654,g26098);
	nor 	XG13697 	(g28353,g24732,g27654,g9073);
	or 	XG13698 	(g28513,g26123,g27276);
	and 	XG13699 	(g26838,g24515,g2860);
	or 	XG13700 	(g29294,g18779,g28645);
	or 	XG13701 	(g28526,g26178,g27285);
	or 	XG13702 	(g28051,g18166,g27699);
	and 	XG13703 	(g25850,g24636,g3502);
	and 	XG13704 	(g27957,g15995,g25947);
	and 	XG13705 	(g27932,g19369,g25944);
	or 	XG13706 	(g29271,g18637,g28333);
	or 	XG13707 	(g29305,g18811,g28602);
	or 	XG13708 	(g29261,g18605,g28247);
	and 	XG13709 	(g26839,g24516,g2988);
	or 	XG13710 	(g29308,g18815,g28612);
	and 	XG13711 	(g28152,g27279,g26297);
	or 	XG13712 	(g28561,g26250,g27312);
	or 	XG13713 	(g28594,g26289,g27334);
	or 	XG13714 	(g28525,g26176,g27284);
	or 	XG13715 	(g29267,g18622,g28257);
	not 	XG13716 	(g26818,I25530);
	not 	XG13717 	(g29190,g27046);
	or 	XG13718 	(g29288,g18762,g28630);
	and 	XG13719 	(g26847,g24525,g2873);
	or 	XG13720 	(g28546,g26231,g27302);
	or 	XG13721 	(g28058,g18268,g27235);
	or 	XG13722 	(g28607,g26303,g27342);
	or 	XG13723 	(g28596,g26291,g27336);
	and 	XG13724 	(g26287,g25225,g2138);
	and 	XG13725 	(g26279,g25213,g4249);
	or 	XG13726 	(g28517,g26154,g27280);
	and 	XG13727 	(g26846,g24524,g37);
	or 	XG13728 	(g28565,g26253,g27315);
	or 	XG13729 	(g29290,g18764,g28569);
	or 	XG13730 	(g29287,g18760,g28555);
	or 	XG13731 	(g28566,g26254,g27316);
	and 	XG13732 	(g26854,g24534,g2868);
	and 	XG13733 	(g26294,g25230,g4245);
	or 	XG13734 	(g28047,g18160,g27676);
	and 	XG13735 	(g26292,g25228,g2689);
	or 	XG13736 	(g28560,g26249,g27311);
	or 	XG13737 	(g29289,g18763,g28642);
	or 	XG13738 	(g29281,g18743,g28541);
	and 	XG13739 	(g26849,g24527,g2994);
	or 	XG13740 	(g28050,g18165,g27692);
	or 	XG13741 	(g28049,g18164,g27684);
	and 	XG13742 	(g26848,g24526,g2950);
	or 	XG13743 	(g28046,g18157,g27667);
	or 	XG13744 	(g28562,g26251,g27313);
	or 	XG13745 	(g28589,g26285,g27331);
	and 	XG13746 	(g26304,g25246,g2697);
	and 	XG13747 	(g25782,g24571,g2936);
	and 	XG13748 	(g25775,g24568,g2922);
	and 	XG13749 	(g26853,g24533,g94);
	or 	XG13750 	(g29260,g18604,g28315);
	and 	XG13751 	(g26312,g25264,g2704);
	and 	XG13752 	(g25768,g24560,g2912);
	not 	XG13753 	(g28479,g27654);
	and 	XG13754 	(g26257,g25197,g4253);
	or 	XG13755 	(g29259,g18603,g28304);
	and 	XG13756 	(g26842,g24522,g2894);
	or 	XG13757 	(g28625,g26324,g27363);
	or 	XG13758 	(g29258,g18601,g28238);
	or 	XG13759 	(g28614,g26311,g27351);
	and 	XG13760 	(g26858,g24540,g2970);
	or 	XG13761 	(g27224,g15678,g25870);
	nand 	XG13762 	(I24363,g14320,g23687);
	and 	XG13763 	(g28198,g27492,g26649);
	or 	XG13764 	(g27250,g15738,g25901);
	or 	XG13765 	(g27016,g14585,g26821);
	and 	XG13766 	(g27393,g20066,g26099);
	or 	XG13767 	(g29643,g27145,g28192);
	and 	XG13768 	(g27964,g22492,g25956);
	and 	XG13769 	(g27968,g19614,g25958);
	and 	XG13770 	(g27612,g8844,g25887);
	or 	XG13771 	(g28533,g26203,g27291);
	nor 	XG13772 	(g29933,g12259,g28500,g8808);
	and 	XG13773 	(g29475,g28500,g14033);
	nand 	XG13774 	(I22923,I22921,g21284);
	and 	XG13775 	(g24949,g20751,g23796);
	or 	XG13776 	(g27024,g17692,g26826);
	and 	XG13777 	(g28573,g27059,g7349);
	nand 	XG13778 	(g28174,g27059,g1270);
	and 	XG13779 	(g28653,g27014,g7544);
	or 	XG13780 	(g28538,g26206,g27294);
	and 	XG13781 	(g24912,g20682,g23687);
	and 	XG13782 	(g28160,g27463,g26309);
	not 	XG13783 	(g28325,g27463);
	nand 	XG13784 	(I24461,g14437,g23796);
	not 	XG13785 	(g30184,g28144);
	and 	XG13786 	(g24939,g21012,g23771);
	nand 	XG13787 	(I23978,g13670,g23198);
	not 	XG13788 	(g29196,g27059);
	and 	XG13789 	(g28597,g20508,g27515);
	not 	XG13790 	(I26989,g27277);
	or 	XG13791 	(g28527,g26182,g27286);
	or 	XG13792 	(g27026,g17726,g26828);
	not 	XG13793 	(g28431,I26925);
	and 	XG13794 	(g28164,g27528,g8651);
	nand 	XG13795 	(g28504,g11679,g27528,g758);
	nand 	XG13796 	(I23917,g9333,g23975);
	or 	XG13797 	(g29325,g27820,g28813);
	or 	XG13798 	(g28279,g25909,g27087);
	nand 	XG13799 	(I24438,g14411,g23771);
	not 	XG13800 	(g29745,g28500);
	or 	XG13801 	(g28368,g27184,g27158);
	not 	XG13802 	(g28370,g27528);
	and 	XG13803 	(g27036,g11038,g26329);
	and 	XG13804 	(g27043,g8632,g26335);
	and 	XG13805 	(g27035,g1500,g26348);
	and 	XG13806 	(g27030,g7947,g26343);
	and 	XG13807 	(g24564,g21163,g23198);
	nor 	XG13808 	(g28444,g24825,g27463,g8575);
	and 	XG13809 	(g29477,g28441,g14090);
	or 	XG13810 	(g27231,g15699,g25873);
	or 	XG13811 	(g27258,g15749,g25905);
	or 	XG13812 	(g29319,g14453,g28812);
	and 	XG13813 	(g30173,g13082,g28118);
	and 	XG13814 	(g28314,g14205,g27552);
	and 	XG13815 	(g28285,g27717,g9657);
	and 	XG13816 	(g28672,g27017,g7577);
	not 	XG13817 	(g28598,g27717);
	or 	XG13818 	(g29114,g26602,g27646);
	and 	XG13819 	(g28237,g27597,g9492);
	not 	XG13820 	(g25838,g25250);
	not 	XG13821 	(I25562,g25250);
	not 	XG13822 	(g25783,g25250);
	not 	XG13823 	(g25869,g25250);
	or 	XG13824 	(g28180,g27511,g20242);
	not 	XG13825 	(I26710,g27511);
	not 	XG13826 	(I27492,g27511);
	not 	XG13827 	(g28119,g27008);
	nand 	XG13828 	(I25221,I25219,g24718);
	not 	XG13829 	(g26827,g24819);
	not 	XG13830 	(g26831,g24836);
	not 	XG13831 	(g26832,g24850);
	not 	XG13832 	(g26837,g24869);
	not 	XG13833 	(g25790,g25027);
	not 	XG13834 	(g25820,g25051);
	not 	XG13835 	(I25146,g24911);
	not 	XG13836 	(I25161,g24920);
	not 	XG13837 	(g25837,g25064);
	not 	XG13838 	(g26836,g24866);
	not 	XG13839 	(g26841,g24893);
	nand 	XG13840 	(I25244,I25242,g24744);
	or 	XG13841 	(g26082,g24561,g2898);
	not 	XG13842 	(g26364,I25327);
	not 	XG13843 	(I24759,g24229);
	not 	XG13844 	(I24839,g24298);
	not 	XG13845 	(I25677,g25640);
	nand 	XG13846 	(I25220,I25219,g482);
	not 	XG13847 	(g26483,I25359);
	or 	XG13848 	(g26874,I25613,I25612);
	or 	XG13849 	(g26365,g25141,g25504);
	not 	XG13850 	(g24891,g23231);
	nor 	XG13851 	(g27366,g26636,g8016);
	and 	XG13852 	(g26604,g25051,g13248);
	and 	XG13853 	(g26547,g25027,g13283);
	nor 	XG13854 	(g27027,g26484,g26398);
	nor 	XG13855 	(g26976,g25791,g5016);
	nor 	XG13856 	(g27400,g26657,g8553);
	and 	XG13857 	(g26541,g24375,g319);
	nor 	XG13858 	(g27703,g25791,g9607);
	nor 	XG13859 	(g27771,g25839,g9809);
	nor 	XG13860 	(g27368,g26657,g8119);
	and 	XG13861 	(g26381,g25548,g4456);
	not 	XG13862 	(g25240,g23650);
	nor 	XG13863 	(g27875,g25821,g9875);
	nor 	XG13864 	(g27954,g25856,g10014);
	nor 	XG13865 	(g27770,g25821,g9386);
	nor 	XG13866 	(g27823,g25805,g9792);
	and 	XG13867 	(g25765,g24973,g24989);
	nand 	XG13868 	(g28796,g7335,g7418,g27858);
	nand 	XG13869 	(g28966,g7380,g2361,g27858);
	nor 	XG13870 	(g27704,g25791,g7239);
	nor 	XG13871 	(g27354,g26636,g8064);
	or 	XG13872 	(g25774,g12043,g25223);
	and 	XG13873 	(g26511,g24364,g19265);
	nor 	XG13874 	(g27926,g25856,g9467);
	nand 	XG13875 	(g24808,I23987,I23986);
	nand 	XG13876 	(g28843,g7387,g7456,g27907);
	nand 	XG13877 	(g28874,g2421,g7424,g27907);
	nand 	XG13878 	(g28837,g2197,g7374,g27800);
	nand 	XG13879 	(g28903,g7280,g2197,g27800);
	nor 	XG13880 	(g27722,g25805,g7247);
	not 	XG13881 	(g25260,I24448);
	nor 	XG13882 	(g27927,g25856,g9621);
	or 	XG13883 	(g29248,g18434,g28677);
	and 	XG13884 	(g25780,g25527,g25532);
	nand 	XG13885 	(g24380,I23602,I23601);
	and 	XG13886 	(g26166,g7558,g11709,g11724,g25357);
	and 	XG13887 	(g26148,g11686,g11709,g11724,g25357);
	not 	XG13888 	(g25180,g23529);
	nor 	XG13889 	(g27382,g26657,g8219);
	not 	XG13890 	(g25380,g23776);
	and 	XG13891 	(g26819,g24490,g106);
	nor 	XG13892 	(g27982,g25856,g7212);
	nand 	XG13893 	(g28765,g7280,g7374,g27800);
	nand 	XG13894 	(g28935,g7328,g2227,g27800);
	not 	XG13895 	(g25296,g23745);
	not 	XG13896 	(g26860,I25594);
	not 	XG13897 	(g25241,g23651);
	and 	XG13898 	(g26190,g11686,g7586,g11724,g25357);
	and 	XG13899 	(g26213,g7558,g7586,g11724,g25357);
	and 	XG13900 	(g26308,g25289,g6961);
	nor 	XG13901 	(g27826,g25821,g9501);
	and 	XG13902 	(g26630,g24419,g7592);
	and 	XG13903 	(g26652,g24426,g10799);
	nand 	XG13904 	(g28871,g2331,g7418,g27858);
	nand 	XG13905 	(g28942,g7335,g2331,g27858);
	and 	XG13906 	(g26358,g25528,g19522);
	and 	XG13907 	(g26394,g25560,g22530);
	and 	XG13908 	(g26399,g25566,g15572);
	nor 	XG13909 	(g27924,g25839,g9946);
	not 	XG13910 	(g24759,g23003);
	and 	XG13911 	(g26380,g25547,g19572);
	and 	XG13912 	(g26379,g25546,g19904);
	and 	XG13913 	(g26357,g25525,g22547);
	and 	XG13914 	(g26395,g25561,g22547);
	and 	XG13915 	(g26391,g25555,g19593);
	and 	XG13916 	(g26389,g25553,g19949);
	nor 	XG13917 	(g27647,g26616,g3004);
	and 	XG13918 	(g26857,g25049,g25062);
	nor 	XG13919 	(g27828,g25856,g9892);
	not 	XG13920 	(g24417,g22171);
	nor 	XG13921 	(g27829,g25856,g7345);
	and 	XG13922 	(g26612,g24407,g901);
	nand 	XG13923 	(g28946,g2421,g2495,g27907);
	nand 	XG13924 	(g28994,g7424,g2495,g27907);
	nand 	XG13925 	(g29131,g9762,g27907);
	nand 	XG13926 	(g29134,g27907,g9762);
	not 	XG13927 	(g26856,I25586);
	and 	XG13928 	(g26852,g24958,g24975);
	or 	XG13929 	(g29225,g18158,g28451);
	not 	XG13930 	(g25298,g23760);
	and 	XG13931 	(g26871,g25020,g25038);
	nor 	XG13932 	(g27010,g25839,g6052);
	nor 	XG13933 	(g27879,g25856,g9523);
	not 	XG13934 	(I26667,g27585);
	and 	XG13935 	(g25772,g24934,g24944);
	nor 	XG13936 	(g27337,g26616,g8334);
	not 	XG13937 	(g23684,I22819);
	and 	XG13938 	(g28236,g27971,g8515);
	and 	XG13939 	(g28245,g27975,g11367);
	nor 	XG13940 	(g27721,g25805,g9672);
	and 	XG13941 	(g26863,g24957,g24974);
	or 	XG13942 	(g25767,g12015,g25207);
	nand 	XG13943 	(g28867,g2153,g2227,g27800);
	nand 	XG13944 	(g28793,g2153,g7328,g27800);
	nand 	XG13945 	(g29057,g9649,g27800);
	nand 	XG13946 	(g29060,g27800,g9649);
	nand 	XG13947 	(I25908,I25907,g26256);
	nand 	XG13948 	(I25909,I25907,g24782);
	and 	XG13949 	(g26513,g24365,g19501);
	and 	XG13950 	(g26650,g24424,g10796);
	and 	XG13951 	(g26542,g24376,g13102);
	and 	XG13952 	(g26651,g24425,g22707);
	and 	XG13953 	(g26670,g24428,g13385);
	and 	XG13954 	(g26671,g24429,g316);
	and 	XG13955 	(g27599,g20033,g26337);
	and 	XG13956 	(I26960,g22698,g26424,g24995);
	and 	XG13957 	(I27409,g22698,g26424,g25556);
	and 	XG13958 	(I27381,g22698,g26424,g25549);
	and 	XG13959 	(I27429,g22698,g26424,g25562);
	and 	XG13960 	(I27364,g22698,g26424,g25541);
	and 	XG13961 	(I26972,g22698,g26424,g25011);
	and 	XG13962 	(I27349,g22698,g26424,g25534);
	and 	XG13963 	(I26948,g22698,g26424,g24981);
	nor 	XG13964 	(g27356,g26657,g9429);
	nor 	XG13965 	(g27338,g26616,g9291);
	and 	XG13966 	(g26689,g24431,g15754);
	and 	XG13967 	(g26360,g25533,g10589);
	nor 	XG13968 	(g27732,g25791,g9364);
	and 	XG13969 	(g26517,g24367,g15708);
	nor 	XG13970 	(g27735,g25821,g7262);
	nand 	XG13971 	(I25846,I25845,g26212);
	nand 	XG13972 	(I25847,I25845,g24799);
	and 	XG13973 	(g26571,g24386,g10472);
	and 	XG13974 	(g26543,g24377,g12910);
	nor 	XG13975 	(g27733,g25805,g9305);
	and 	XG13976 	(g26486,g24358,g4423);
	and 	XG13977 	(g26390,g25554,g4423);
	not 	XG13978 	(g25272,g23715);
	and 	XG13979 	(g26393,g25558,g19467);
	and 	XG13980 	(g26347,g24850,g262);
	nor 	XG13981 	(g27768,g25805,g9264);
	nor 	XG13982 	(g27364,g26616,g8426);
	and 	XG13983 	(g26258,g25231,g12875);
	and 	XG13984 	(g26356,g25523,g15581);
	and 	XG13985 	(g26325,g25370,g12644);
	nor 	XG13986 	(g27343,g26616,g8005);
	and 	XG13987 	(g26613,g24518,g1361);
	or 	XG13988 	(g25917,g24518,g22524);
	not 	XG13989 	(g25221,g23653);
	and 	XG13990 	(g26362,g25538,g19557);
	and 	XG13991 	(g26378,g25544,g19576);
	nor 	XG13992 	(g27966,g25805,g7153);
	and 	XG13993 	(g26200,g10627,g10658,g10678,g24688);
	and 	XG13994 	(g26241,g10627,g8778,g10678,g24688);
	and 	XG13995 	(g26313,g25326,g12645);
	and 	XG13996 	(g26423,g24356,g19488);
	not 	XG13997 	(I25692,g25689);
	nor 	XG13998 	(g27353,g26616,g8097);
	nor 	XG13999 	(g27659,g26657,g3706);
	not 	XG14000 	(g25781,g24510);
	and 	XG14001 	(g26861,g25003,g25021);
	nor 	XG14002 	(g27731,g25791,g9229);
	and 	XG14003 	(g26388,g25552,g19595);
	not 	XG14004 	(g25206,g23613);
	not 	XG14005 	(g25513,g23870);
	nor 	XG14006 	(g27516,g26657,g9180);
	not 	XG14007 	(I24278,g23440);
	not 	XG14008 	(I24281,g23440);
	not 	XG14009 	(I25683,g25642);
	not 	XG14010 	(I25695,g25690);
	nor 	XG14011 	(g27960,g25791,g7134);
	nor 	XG14012 	(g27007,g25821,g5706);
	and 	XG14013 	(g26261,g8757,g8778,g10678,g24688);
	and 	XG14014 	(g26223,g8757,g10658,g10678,g24688);
	not 	XG14015 	(g25786,g24518);
	nor 	XG14016 	(g27969,g25821,g7170);
	nor 	XG14017 	(g27720,g25791,g9253);
	and 	XG14018 	(g26339,g24836,g225);
	and 	XG14019 	(g26397,g25563,g19475);
	and 	XG14020 	(g26487,g24359,g15702);
	not 	XG14021 	(g29170,g27907);
	not 	XG14022 	(g29152,g27907);
	not 	XG14023 	(g29130,g27907);
	not 	XG14024 	(g28713,g27907);
	and 	XG14025 	(g26351,g24869,g239);
	not 	XG14026 	(g25297,g23746);
	and 	XG14027 	(g26244,g8757,g10658,g8812,g24688);
	and 	XG14028 	(g26281,g8757,g8778,g8812,g24688);
	and 	XG14029 	(g26226,g10627,g10658,g8812,g24688);
	and 	XG14030 	(g26264,g10627,g8778,g8812,g24688);
	and 	XG14031 	(g26753,g24452,g16024);
	and 	XG14032 	(g26719,g24438,g10709);
	and 	XG14033 	(g26336,g25480,g10307);
	nand 	XG14034 	(g28907,g2287,g2361,g27858);
	nand 	XG14035 	(g28840,g2287,g7380,g27858);
	nand 	XG14036 	(g29097,g27858,g9700);
	nand 	XG14037 	(g29094,g9700,g27858);
	not 	XG14038 	(g29092,g27800);
	not 	XG14039 	(g29056,g27800);
	not 	XG14040 	(g29128,g27800);
	not 	XG14041 	(g28678,g27800);
	not 	XG14042 	(g28696,g27858);
	not 	XG14043 	(g29093,g27858);
	not 	XG14044 	(g29129,g27858);
	not 	XG14045 	(g29151,g27858);
	not 	XG14046 	(g23453,I22576);
	not 	XG14047 	(g25424,g23800);
	not 	XG14048 	(I25680,g25641);
	not 	XG14049 	(g25465,g23824);
	nand 	XG14050 	(g24369,I23587,I23586);
	or 	XG14051 	(g29227,g18169,g28456);
	and 	XG14052 	(g26259,g25232,g24430);
	and 	XG14053 	(g27369,g25324,g25894);
	not 	XG14054 	(I24237,g23823);
	nand 	XG14055 	(I25243,I25242,g490);
	nand 	XG14056 	(g24802,I23971,I23970);
	not 	XG14057 	(I25786,g26424);
	not 	XG14058 	(I25779,g26424);
	not 	XG14059 	(I25790,g26424);
	not 	XG14060 	(g27730,g26424);
	not 	XG14061 	(I25689,g25688);
	and 	XG14062 	(g26306,g25286,g13087);
	and 	XG14063 	(g26350,g25517,g13087);
	and 	XG14064 	(g26295,g25266,g13070);
	and 	XG14065 	(g26307,g25288,g13070);
	and 	XG14066 	(g26345,g25505,g13051);
	and 	XG14067 	(g26280,g25248,g13051);
	and 	XG14068 	(g26610,g24405,g14198);
	and 	XG14069 	(g26629,g24418,g14173);
	and 	XG14070 	(g27697,g23649,g25785);
	and 	XG14071 	(g27696,g23647,g25800);
	and 	XG14072 	(g30125,g21056,g28581);
	and 	XG14073 	(g27673,g23541,g25769);
	and 	XG14074 	(g27674,g23543,g26873);
	and 	XG14075 	(g27288,g23013,g26515);
	and 	XG14076 	(g27287,g23011,g26545);
	and 	XG14077 	(g30110,g20916,g28564);
	and 	XG14078 	(g30135,g21180,g28592);
	and 	XG14079 	(g30066,g20636,g28518);
	and 	XG14080 	(g30099,g20776,g28549);
	and 	XG14081 	(g27683,g23567,g25770);
	and 	XG14082 	(g27682,g23565,g25777);
	and 	XG14083 	(g28178,g19397,g27019);
	and 	XG14084 	(g27665,g23519,g26872);
	and 	XG14085 	(g27666,g23521,g26865);
	and 	XG14086 	(g30094,g20767,g28544);
	and 	XG14087 	(g30084,g20700,g28534);
	and 	XG14088 	(g27299,g23028,g26546);
	and 	XG14089 	(g27298,g23026,g26573);
	and 	XG14090 	(g30095,g20768,g28545);
	and 	XG14091 	(g27691,g23609,g25778);
	and 	XG14092 	(g27690,g23607,g25784);
	and 	XG14093 	(g27310,g23059,g26574);
	and 	XG14094 	(g27309,g23057,g26603);
	and 	XG14095 	(g30121,g21052,g28577);
	and 	XG14096 	(g30086,g20704,g28536);
	and 	XG14097 	(g30122,g21054,g28578);
	and 	XG14098 	(g30133,g21179,g28591);
	and 	XG14099 	(g30158,g21274,g28613);
	and 	XG14100 	(g27660,g22763,g26424,g24688);
	nor 	XG14101 	(g27766,g25791,g9716);
	nor 	XG14102 	(g27479,g26616,g9056);
	nand 	XG14103 	(g29049,g27779,g9640);
	nand 	XG14104 	(g29046,g9640,g27779);
	nand 	XG14105 	(g28857,g1728,g1802,g27779);
	nand 	XG14106 	(g28920,g7315,g1802,g27779);
	nor 	XG14107 	(g27652,g26636,g3355);
	nor 	XG14108 	(g27827,g25839,g9456);
	nor 	XG14109 	(g27772,g25839,g7297);
	nand 	XG14110 	(I23950,I23949,g23162);
	nor 	XG14111 	(g27877,g25839,g9397);
	nor 	XG14112 	(g27973,g25839,g7187);
	nor 	XG14113 	(g27367,g26636,g8155);
	or 	XG14114 	(g29275,g21868,g28165);
	nand 	XG14115 	(I24384,I24383,g23721);
	nor 	XG14116 	(g27352,g26616,g7975);
	nor 	XG14117 	(g26993,g25805,g5360);
	nor 	XG14118 	(g27345,g26636,g9360);
	nor 	XG14119 	(g27012,g25856,g6398);
	or 	XG14120 	(g26800,g24929,g24922);
	nor 	XG14121 	(g27734,g25821,g9733);
	nand 	XG14122 	(g28911,g2465,g7456,g27907);
	nand 	XG14123 	(g28973,g7387,g2465,g27907);
	nand 	XG14124 	(g28783,g1728,g7315,g27779);
	nand 	XG14125 	(g28758,g7275,g7356,g27779);
	nand 	XG14126 	(I24415,I24414,g23751);
	nor 	XG14127 	(g27825,g25821,g9316);
	nand 	XG14128 	(g25996,g22838,g24601);
	nor 	XG14129 	(g27355,g26657,g8443);
	and 	XG14130 	(g28547,g27091,g6821);
	and 	XG14131 	(g28524,g27084,g6821);
	and 	XG14132 	(g28535,g27088,g11981);
	and 	XG14133 	(g28563,g27100,g11981);
	nor 	XG14134 	(g27381,g26657,g8075);
	and 	XG14135 	(g28537,g27089,g6832);
	and 	XG14136 	(g28567,g27101,g6832);
	and 	XG14137 	(g28550,g27092,g12009);
	and 	XG14138 	(g28583,g27112,g12009);
	or 	XG14139 	(g25911,g24510,g22514);
	and 	XG14140 	(g26606,g24510,g1018);
	and 	XG14141 	(g26236,g7558,g7586,g6856,g25357);
	and 	XG14142 	(g26218,g11686,g7586,g6856,g25357);
	and 	XG14143 	(g26195,g7558,g11709,g6856,g25357);
	and 	XG14144 	(g26171,g11686,g11709,g6856,g25357);
	nand 	XG14145 	(I24416,I24414,g14382);
	and 	XG14146 	(g28268,g27990,g8572);
	and 	XG14147 	(g28246,g27976,g8572);
	and 	XG14148 	(g28284,g27994,g11398);
	and 	XG14149 	(g28256,g27984,g11398);
	nand 	XG14150 	(g28824,g1772,g7356,g27779);
	nand 	XG14151 	(g28892,g7275,g1772,g27779);
	nor 	XG14152 	(g27769,g25805,g9434);
	nor 	XG14153 	(g27344,g26636,g8390);
	not 	XG14154 	(g29115,g27779);
	not 	XG14155 	(g29080,g27779);
	not 	XG14156 	(g29045,g27779);
	not 	XG14157 	(g28675,g27779);
	not 	XG14158 	(g26187,I25190);
	not 	XG14159 	(g28656,g27742);
	not 	XG14160 	(g29079,g27742);
	not 	XG14161 	(g29014,g27742);
	not 	XG14162 	(g29044,g27742);
	or 	XG14163 	(g28208,g27028,g27025);
	nor 	XG14164 	(g27379,g26636,g8492);
	nor 	XG14165 	(g27878,g25839,g9559);
	not 	XG14166 	(g28121,g27093);
	not 	XG14167 	(g28127,g27102);
	nor 	XG14168 	(g27499,g26636,g9095);
	not 	XG14169 	(g25168,I24334);
	not 	XG14170 	(I26654,g27576);
	or 	XG14171 	(g28134,g27962,g27958);
	nand 	XG14172 	(I24385,I24383,g14347);
	nor 	XG14173 	(g28149,g27612,g27598);
	not 	XG14174 	(I27192,g27662);
	or 	XG14175 	(g24952,I24117,g21340,g21326);
	nor 	XG14176 	(g27063,g26516,g26485);
	not 	XG14177 	(g24483,I23688);
	not 	XG14178 	(g25284,I24474);
	not 	XG14179 	(g24489,I23694);
	not 	XG14180 	(g24481,I23684);
	not 	XG14181 	(g24477,I23680);
	not 	XG14182 	(g25265,I24455);
	not 	XG14183 	(g24466,I23671);
	not 	XG14184 	(g25322,I24497);
	not 	XG14185 	(g26326,g24872);
	not 	XG14186 	(g25849,g24491);
	not 	XG14187 	(g25893,g24541);
	not 	XG14188 	(g25886,g24537);
	not 	XG14189 	(g25830,g24485);
	nand 	XG14190 	(g28830,g7369,g7451,g27886);
	nand 	XG14191 	(g28864,g1996,g7411,g27886);
	or 	XG14192 	(g29242,g18354,g28674);
	nand 	XG14193 	(I23951,I23949,g13603);
	nand 	XG14194 	(g25984,g22668,g24567);
	or 	XG14195 	(g29247,g18410,g28694);
	or 	XG14196 	(g29246,g18406,g28710);
	nand 	XG14197 	(g25995,g22853,g24621);
	or 	XG14198 	(g29230,g18202,g28107);
	or 	XG14199 	(g26781,g24921,g24913);
	or 	XG14200 	(g29243,g18358,g28657);
	or 	XG14201 	(g29223,g18131,g28341);
	nand 	XG14202 	(g28853,g7252,g1636,g27742);
	nand 	XG14203 	(g28780,g1636,g7308,g27742);
	or 	XG14204 	(g29255,g18516,g28714);
	or 	XG14205 	(g29241,g18332,g28638);
	nand 	XG14206 	(g28736,g7252,g7308,g27742);
	nand 	XG14207 	(g28755,g1592,g7268,g27742);
	or 	XG14208 	(g28048,g18163,g27362);
	nand 	XG14209 	(g28931,g1996,g2070,g27886);
	nand 	XG14210 	(g28987,g7411,g2070,g27886);
	nand 	XG14211 	(g29118,g9755,g27886);
	nand 	XG14212 	(g29121,g27886,g9755);
	or 	XG14213 	(g29253,g18490,g28697);
	nand 	XG14214 	(g23778,I22923,I22922);
	or 	XG14215 	(g29226,g18159,g28455);
	or 	XG14216 	(g29235,g18260,g28110);
	and 	XG14217 	(g30049,g28167,g13114);
	nor 	XG14218 	(g29359,g28167,g7528);
	and 	XG14219 	(g28255,g27983,g8515);
	and 	XG14220 	(g28265,g27989,g11367);
	or 	XG14221 	(g29240,g18328,g28655);
	not 	XG14222 	(I26004,g26818);
	or 	XG14223 	(g29245,g18384,g28676);
	nand 	XG14224 	(g28927,g7322,g1906,g27837);
	nand 	XG14225 	(g28861,g1906,g7405,g27837);
	nand 	XG14226 	(g28877,g7431,g7490,g27937);
	nand 	XG14227 	(g28914,g2555,g7462,g27937);
	or 	XG14228 	(g29229,g18191,g28532);
	or 	XG14229 	(g26278,g24549,g24545);
	or 	XG14230 	(g29250,g18460,g28695);
	or 	XG14231 	(g28132,g27957,g27932);
	nand 	XG14232 	(g28900,g2040,g7451,g27886);
	nand 	XG14233 	(g28962,g7369,g2040,g27886);
	nand 	XG14234 	(g29660,g9582,g28448);
	nand 	XG14235 	(g28885,g7268,g1668,g27742);
	nand 	XG14236 	(g28820,g1592,g1668,g27742);
	nand 	XG14237 	(g29015,g9586,g27742);
	nand 	XG14238 	(g29018,g27742,g9586);
	nand 	XG14239 	(g28786,g7322,g7405,g27837);
	nand 	XG14240 	(g28955,g7362,g1936,g27837);
	or 	XG14241 	(g24240,g18251,g22861);
	not 	XG14242 	(g29507,g28353);
	or 	XG14243 	(g29254,g18512,g28725);
	or 	XG14244 	(g30334,g18143,g29837);
	nand 	XG14245 	(g25985,g23956,g24631);
	nand 	XG14246 	(g26025,g24631,g22405);
	nand 	XG14247 	(g25953,g22688,g24570,g22756);
	nand 	XG14248 	(g26052,g22921,g24662,g22714);
	or 	XG14249 	(g26293,g24555,g24550);
	or 	XG14250 	(g24241,g18252,g22920);
	nand 	XG14251 	(g29025,g7462,g2629,g27937);
	nand 	XG14252 	(g28977,g2555,g2629,g27937);
	nand 	XG14253 	(g29154,g9835,g27937);
	nand 	XG14254 	(g29157,g27937,g9835);
	and 	XG14255 	(g30671,g22317,g29319);
	and 	XG14256 	(g29378,g22493,g28137);
	or 	XG14257 	(g24257,g18310,g22938);
	or 	XG14258 	(g29251,g18464,g28679);
	nand 	XG14259 	(g29001,g7431,g2599,g27937);
	nand 	XG14260 	(g28950,g2599,g7490,g27937);
	not 	XG14261 	(g29177,g27937);
	not 	XG14262 	(g29171,g27937);
	not 	XG14263 	(g28726,g27937);
	not 	XG14264 	(g29153,g27937);
	nand 	XG14265 	(I23962,I23961,g23184);
	not 	XG14266 	(g29149,g27837);
	not 	XG14267 	(g29081,g27837);
	not 	XG14268 	(g29116,g27837);
	not 	XG14269 	(g28693,g27837);
	not 	XG14270 	(g28711,g27886);
	not 	XG14271 	(g29117,g27886);
	not 	XG14272 	(g29169,g27886);
	not 	XG14273 	(g29150,g27886);
	and 	XG14274 	(g29513,g14095,g28448);
	or 	XG14275 	(g29228,g18173,g28426);
	or 	XG14276 	(g28211,g27034,g27029);
	not 	XG14277 	(g29333,g28167);
	or 	XG14278 	(g29252,g18486,g28712);
	or 	XG14279 	(g29244,g18380,g28692);
	and 	XG14280 	(g29834,g23278,g28368);
	or 	XG14281 	(g24256,g18309,g22873);
	or 	XG14282 	(g28135,g27963,g27959);
	nand 	XG14283 	(I23963,I23961,g13631);
	or 	XG14284 	(g29249,g18438,g28658);
	or 	XG14285 	(g29583,g27099,g28182);
	and 	XG14286 	(g30089,g20709,g28538);
	and 	XG14287 	(g30126,g21058,g28582);
	and 	XG14288 	(g30137,g21181,g28594);
	and 	XG14289 	(g30161,g21275,g28614);
	and 	XG14290 	(g28442,g20072,g27278);
	and 	XG14291 	(g28626,g20573,g27542);
	and 	XG14292 	(g30078,g20667,g28526);
	and 	XG14293 	(g30112,g20919,g28566);
	and 	XG14294 	(g30124,g21055,g28580);
	and 	XG14295 	(g30149,g21248,g28605);
	and 	XG14296 	(g30111,g20917,g28565);
	and 	XG14297 	(g30098,g20774,g28548);
	and 	XG14298 	(g28185,g19435,g27026);
	and 	XG14299 	(g28440,g20059,g27274);
	and 	XG14300 	(g28616,g20551,g27532);
	and 	XG14301 	(g30109,g20912,g28562);
	and 	XG14302 	(g30075,g20662,g28525);
	and 	XG14303 	(g30145,g21247,g28603);
	and 	XG14304 	(g30120,g21051,g28576);
	and 	XG14305 	(g30108,g20910,g28561);
	and 	XG14306 	(g30051,g20604,g28513);
	and 	XG14307 	(g30083,g20698,g28533);
	and 	XG14308 	(g30118,g21050,g28574);
	and 	XG14309 	(g28301,g19750,g27224);
	and 	XG14310 	(g28415,g19963,g27250);
	and 	XG14311 	(g28183,g19421,g27024);
	and 	XG14312 	(g28171,g19385,g27016);
	and 	XG14313 	(g29324,g18883,g29078);
	and 	XG14314 	(g30107,g20909,g28560);
	and 	XG14315 	(g30064,g20630,g28517);
	and 	XG14316 	(g30131,g21178,g28589);
	and 	XG14317 	(g30096,g20770,g28546);
	and 	XG14318 	(g30139,g21184,g28596);
	and 	XG14319 	(g30101,g20780,g28551);
	and 	XG14320 	(g30172,g21286,g28625);
	and 	XG14321 	(g30151,g21249,g28607);
	and 	XG14322 	(g30138,g21182,g28595);
	and 	XG14323 	(g31252,g20101,g29643);
	and 	XG14324 	(g29746,g20037,g28279);
	nand 	XG14325 	(g25974,g22837,g24576);
	nand 	XG14326 	(I24439,I24438,g23771);
	and 	XG14327 	(g29367,g28325,g8575);
	nand 	XG14328 	(g29082,g9694,g27837);
	nand 	XG14329 	(g29085,g27837,g9694);
	nand 	XG14330 	(g28896,g1862,g1936,g27837);
	nand 	XG14331 	(g28827,g1862,g7362,g27837);
	or 	XG14332 	(g26751,g24912,g24903);
	and 	XG14333 	(g29924,g29190,g13031);
	nor 	XG14334 	(g29916,g11083,g28504,g8681);
	and 	XG14335 	(g29376,g28504,g14002);
	nand 	XG14336 	(I24440,I24438,g14411);
	nand 	XG14337 	(g26053,g22941,g24677,g22875);
	nand 	XG14338 	(I23918,I23917,g23975);
	or 	XG14339 	(g28053,g18168,g27393);
	nand 	XG14340 	(I23979,I23978,g23198);
	not 	XG14341 	(g29707,g28504);
	nand 	XG14342 	(I24462,I24461,g23796);
	not 	XG14343 	(g30322,g28431);
	not 	XG14344 	(g29744,g28431);
	not 	XG14345 	(I28576,g28431);
	nand 	XG14346 	(g29679,g23042,g28353,g153);
	and 	XG14347 	(g29329,g28353,g7995);
	not 	XG14348 	(g28508,I26989);
	or 	XG14349 	(g29256,g18533,g28597);
	or 	XG14350 	(g26809,g24939,g24930);
	nand 	XG14351 	(I24364,I24363,g23687);
	and 	XG14352 	(g29494,g28479,g9073);
	nand 	XG14353 	(I24463,I24461,g14437);
	or 	XG14354 	(g26813,g24949,g24940);
	or 	XG14355 	(g29508,g27041,g28152);
	or 	XG14356 	(g30287,g27677,g28653);
	nand 	XG14357 	(g31509,g12323,g29933,g599);
	and 	XG14358 	(g30982,g29933,g8895);
	not 	XG14359 	(g29343,g28174);
	not 	XG14360 	(g31243,g29933);
	or 	XG14361 	(g28138,g27968,g27964);
	or 	XG14362 	(g29706,g27208,g28198);
	nand 	XG14363 	(I24365,I24363,g14320);
	and 	XG14364 	(g30062,g28174,g13129);
	nor 	XG14365 	(g29361,g28174,g7553);
	and 	XG14366 	(g30935,g29745,g8808);
	and 	XG14367 	(g29330,g18894,g29114);
	and 	XG14368 	(g29937,g29196,g13044);
	or 	XG14369 	(g26305,g24564,g24556);
	nand 	XG14370 	(I23980,I23978,g13670);
	or 	XG14371 	(g30291,g27685,g28672);
	not 	XG14372 	(I28128,g28314);
	and 	XG14373 	(g29668,g14255,g28527);
	and 	XG14374 	(g31654,g13062,g29325);
	and 	XG14375 	(g29375,g28370,g13946);
	nand 	XG14376 	(I23919,I23917,g9333);
	and 	XG14377 	(g28427,g20008,g27258);
	and 	XG14378 	(g28313,g19766,g27231);
	or 	XG14379 	(g31144,g28193,g29477);
	not 	XG14380 	(g29597,g28444);
	or 	XG14381 	(g28212,g27035,g27030);
	or 	XG14382 	(g28216,g27043,g27036);
	nand 	XG14383 	(g29778,g23204,g28444,g294);
	and 	XG14384 	(g29363,g28444,g8458);
	or 	XG14385 	(g30579,g14571,g30173);
	and 	XG14386 	(g29570,g28598,g2763);
	or 	XG14387 	(g29793,g27247,g28237);
	and 	XG14388 	(I26530,g24098,g24097,g24096,g26365);
	and 	XG14389 	(g27649,g25820,g10820);
	and 	XG14390 	(g27627,g25790,g13266);
	not 	XG14391 	(g28040,g26365);
	not 	XG14392 	(g28034,g26365);
	not 	XG14393 	(g28038,g26365);
	not 	XG14394 	(g28039,g26365);
	not 	XG14395 	(g28032,g26365);
	not 	XG14396 	(I26100,g26365);
	not 	XG14397 	(g28033,g26365);
	not 	XG14398 	(g28036,g26365);
	not 	XG14399 	(g28037,g26365);
	nand 	XG14400 	(g26248,I25221,I25220);
	not 	XG14401 	(g26935,I25677);
	not 	XG14402 	(g25692,I24839);
	not 	XG14403 	(g25620,I24759);
	and 	XG14404 	(g27414,g26827,g255);
	and 	XG14405 	(g27467,g26832,g269);
	and 	XG14406 	(g27439,g26831,g232);
	and 	XG14407 	(g27493,g26837,g246);
	nand 	XG14408 	(g26269,I25244,I25243);
	not 	XG14409 	(g26131,I25161);
	not 	XG14410 	(g26105,I25146);
	not 	XG14411 	(I27758,g28119);
	not 	XG14412 	(g29194,I27492);
	not 	XG14413 	(g28187,I26710);
	not 	XG14414 	(g29385,g28180);
	not 	XG14415 	(g26840,I25562);
	and 	XG14416 	(g27042,g19343,g25774);
	and 	XG14417 	(g27033,g19273,g25767);
	or 	XG14418 	(g26881,g24187,g26629);
	or 	XG14419 	(g26880,g24186,g26610);
	or 	XG14420 	(g26961,g24306,g26280);
	or 	XG14421 	(g26966,g24318,g26345);
	or 	XG14422 	(g26968,g24321,g26307);
	or 	XG14423 	(g26962,g24307,g26295);
	or 	XG14424 	(g26967,g24319,g26350);
	or 	XG14425 	(g26963,g24308,g26306);
	nor 	XG14426 	(g28803,g22763,g27730);
	not 	XG14427 	(g26941,I25689);
	not 	XG14428 	(g27074,I25790);
	not 	XG14429 	(g27051,I25779);
	not 	XG14430 	(g27064,I25786);
	and 	XG14431 	(g29954,g28796,g2299);
	and 	XG14432 	(g28223,g17194,g27338);
	and 	XG14433 	(g27057,g26261,g6227,g6219,g7791);
	nor 	XG14434 	(g26314,g24802,g24808);
	or 	XG14435 	(g26886,g24192,g26651);
	nand 	XG14436 	(g27550,g25772,g24943);
	and 	XG14437 	(g29519,g28840,g2295);
	not 	XG14438 	(g25073,I24237);
	and 	XG14439 	(g27032,g26200,g5188,g5180,g7704);
	or 	XG14440 	(g28082,g24315,g27369);
	or 	XG14441 	(g26964,g24316,g26259);
	and 	XG14442 	(g29628,g28648,g27924);
	not 	XG14443 	(I25606,g25465);
	not 	XG14444 	(g26936,I25680);
	not 	XG14445 	(I25598,g25424);
	not 	XG14446 	(I24393,g23453);
	not 	XG14447 	(I24396,g23453);
	or 	XG14448 	(g26946,g24284,g26389);
	and 	XG14449 	(g27185,g1917,g8302,g26190);
	and 	XG14450 	(g29360,g28294,g27364);
	and 	XG14451 	(g28477,g17676,g27966);
	and 	XG14452 	(g27058,g26264,g3530,g3522,g10323);
	and 	XG14453 	(g29576,g28903,g2177);
	and 	XG14454 	(g28197,g11344,g27647);
	not 	XG14455 	(g30088,g29094);
	not 	XG14456 	(g30020,g29097);
	not 	XG14457 	(g30038,g29097);
	not 	XG14458 	(g30079,g29097);
	not 	XG14459 	(g29913,g28840);
	not 	XG14460 	(g29953,g28907);
	and 	XG14461 	(g28115,g22759,g27354);
	or 	XG14462 	(g26965,g24317,g26336);
	and 	XG14463 	(g28499,g17762,g27982);
	or 	XG14464 	(g26892,g24198,g26719);
	and 	XG14465 	(g29883,g29152,g2465);
	and 	XG14466 	(g27045,g26244,g3179,g3171,g10295);
	and 	XG14467 	(g29968,g28843,g2433);
	or 	XG14468 	(g26893,g24199,g26753);
	and 	XG14469 	(g28010,g25535,g26424,g26223,g23032);
	and 	XG14470 	(g28020,g25542,g26424,g26241,g23032);
	and 	XG14471 	(g27617,g24982,g26424,g26264,g23032);
	and 	XG14472 	(g27602,g24966,g26424,g26244,g23032);
	and 	XG14473 	(g27999,g25529,g26424,g26200,g23032);
	and 	XG14474 	(g26977,g25550,g26424,g26261,g23032);
	and 	XG14475 	(g26994,g25557,g26424,g26226,g23032);
	and 	XG14476 	(g27635,g24996,g26424,g26281,g23032);
	and 	XG14477 	(g29612,g28633,g27875);
	and 	XG14478 	(g28478,g12345,g27007);
	or 	XG14479 	(g26900,g24217,g26819);
	or 	XG14480 	(g26908,g24225,g26358);
	not 	XG14481 	(I25579,g25297);
	or 	XG14482 	(g26906,g24223,g26423);
	and 	XG14483 	(g28454,g12233,g26976);
	or 	XG14484 	(g26956,g24294,g26487);
	nand 	XG14485 	(g27738,g26148,g26424,g25243,g21228);
	nand 	XG14486 	(g27833,g26190,g26424,g25282,g21228);
	nand 	XG14487 	(g27882,g26213,g26424,g25307,g21228);
	nand 	XG14488 	(g27775,g26166,g26424,g25262,g21228);
	or 	XG14489 	(g26905,g24222,g26397);
	and 	XG14490 	(g29364,g28321,g27400);
	or 	XG14491 	(g26902,g24219,g26378);
	and 	XG14492 	(g27044,g26241,g5881,g5873,g7766);
	and 	XG14493 	(g28232,g23586,g27732);
	and 	XG14494 	(g28543,g15628,g27735);
	or 	XG14495 	(g27225,g26364,g2975);
	and 	XG14496 	(g28202,g11413,g27659);
	and 	XG14497 	(g27651,g25781,g22448);
	and 	XG14498 	(g28523,g15585,g27704);
	not 	XG14499 	(g26943,I25695);
	or 	XG14500 	(g26970,g24332,g26308);
	and 	XG14501 	(g29732,g29131,g2514);
	or 	XG14502 	(g30298,g27251,g28245);
	not 	XG14503 	(g26937,I25683);
	not 	XG14504 	(g25115,I24281);
	and 	XG14505 	(g29604,g28966,g2315);
	and 	XG14506 	(g28240,g17239,g27356);
	or 	XG14507 	(g26947,g24285,g26394);
	and 	XG14508 	(g29651,g29134,g2537);
	not 	XG14509 	(I24920,g25513);
	not 	XG14510 	(g26811,g25206);
	or 	XG14511 	(g26952,g24290,g26360);
	or 	XG14512 	(g26903,g24220,g26388);
	or 	XG14513 	(g26904,g24221,g26393);
	or 	XG14514 	(g30293,g27246,g28236);
	and 	XG14515 	(g28272,g26548,g27721);
	and 	XG14516 	(g28139,g26054,g27337);
	not 	XG14517 	(g26942,I25692);
	or 	XG14518 	(g26958,g24297,g26395);
	or 	XG14519 	(g26890,g24196,g26630);
	or 	XG14520 	(g26907,g24224,g26513);
	or 	XG14521 	(g26969,g24329,g26313);
	and 	XG14522 	(g28531,g15608,g27722);
	or 	XG14523 	(g26901,g24218,g26362);
	not 	XG14524 	(g26814,g25221);
	not 	XG14525 	(g27011,g25917);
	and 	XG14526 	(g28116,g26183,g27366);
	nand 	XG14527 	(g27613,g26871,g25048,g24933,g24942);
	or 	XG14528 	(g26971,g24333,g26325);
	or 	XG14529 	(g26945,g24283,g26379);
	or 	XG14530 	(g26949,g24287,g26356);
	or 	XG14531 	(g26960,g24304,g26258);
	and 	XG14532 	(g29588,g28942,g2311);
	and 	XG14533 	(g29596,g28620,g27823);
	or 	XG14534 	(g26889,g24195,g26689);
	not 	XG14535 	(I25567,g25272);
	or 	XG14536 	(g26951,g24289,g26390);
	or 	XG14537 	(g26953,g24291,g26486);
	or 	XG14538 	(g26909,g24227,g26543);
	or 	XG14539 	(g26910,g24228,g26571);
	nand 	XG14540 	(g27141,I25847,I25846);
	and 	XG14541 	(g28225,g23400,g27770);
	or 	XG14542 	(g26954,g24292,g26380);
	or 	XG14543 	(g26957,g24295,g26517);
	or 	XG14544 	(I26522,g26365,g19984,g19935,g19890);
	and 	XG14545 	(g28260,g26518,g27703);
	and 	XG14546 	(g28300,g26605,g27771);
	and 	XG14547 	(g28124,g22842,g27368);
	not 	XG14548 	(I26936,g27599);
	or 	XG14549 	(g26888,g24194,g26671);
	or 	XG14550 	(g26882,g24188,g26650);
	or 	XG14551 	(g26887,g24193,g26542);
	or 	XG14552 	(g26883,g24189,g26670);
	nand 	XG14553 	(g27223,I25909,I25908);
	and 	XG14554 	(g29711,g29134,g2541);
	not 	XG14555 	(g30019,g29060);
	not 	XG14556 	(g30067,g29060);
	not 	XG14557 	(g29997,g29060);
	not 	XG14558 	(g30077,g29057);
	not 	XG14559 	(g29906,g28793);
	not 	XG14560 	(g29942,g28867);
	nand 	XG14561 	(g27931,g25780,g25381,g25425);
	not 	XG14562 	(g25242,g23684);
	and 	XG14563 	(g28489,g12417,g27010);
	not 	XG14564 	(g28156,I26667);
	and 	XG14565 	(g28273,g23729,g27927);
	not 	XG14566 	(g26824,g25298);
	not 	XG14567 	(I26430,g26856);
	not 	XG14568 	(g30039,g29134);
	not 	XG14569 	(g30054,g29134);
	not 	XG14570 	(g30090,g29134);
	not 	XG14571 	(g30100,g29131);
	not 	XG14572 	(g30021,g28994);
	not 	XG14573 	(g29967,g28946);
	and 	XG14574 	(g27759,g26213,g26424,g25224,g22457);
	and 	XG14575 	(g27711,g26166,g26424,g25193,g22369);
	or 	XG14576 	(g27450,g26483,g2917);
	or 	XG14577 	(g26911,g24230,g26612);
	or 	XG14578 	(g26955,g24293,g26391);
	and 	XG14579 	(g29528,g28874,g2429);
	not 	XG14580 	(I25005,g24417);
	and 	XG14581 	(g28244,g26715,g27926);
	nand 	XG14582 	(g27587,g26857,g24918,g25018,g24917);
	and 	XG14583 	(g27724,g26190,g26424,g25208,g22417);
	and 	XG14584 	(g27700,g26148,g26424,g25182,g22342);
	or 	XG14585 	(g26950,g24288,g26357);
	not 	XG14586 	(g26260,g24759);
	or 	XG14587 	(g26948,g24286,g26399);
	not 	XG14588 	(g29981,g28942);
	not 	XG14589 	(g29928,g28871);
	or 	XG14590 	(g26891,g24197,g26652);
	or 	XG14591 	(g27031,g26148,g26166,g26190,g26213);
	and 	XG14592 	(g29525,g28837,g2169);
	not 	XG14593 	(I25555,g25241);
	not 	XG14594 	(I26448,g26860);
	and 	XG14595 	(g27161,g1783,g8241,g26166);
	not 	XG14596 	(I25576,g25296);
	not 	XG14597 	(g29980,g28935);
	not 	XG14598 	(g30299,g28765);
	not 	XG14599 	(I25591,g25380);
	not 	XG14600 	(I25541,g25180);
	and 	XG14601 	(g28599,g8922,g27027);
	not 	XG14602 	(g26816,g25260);
	not 	XG14603 	(g29965,g28903);
	not 	XG14604 	(g29922,g28837);
	not 	XG14605 	(g29923,g28874);
	not 	XG14606 	(g30313,g28843);
	and 	XG14607 	(g29642,g28669,g27954);
	or 	XG14608 	(g26884,g24190,g26511);
	not 	XG14609 	(g29998,g28966);
	not 	XG14610 	(g30306,g28796);
	not 	XG14611 	(I25552,g25240);
	or 	XG14612 	(g26959,g24299,g26381);
	or 	XG14613 	(g26885,g24191,g26541);
	not 	XG14614 	(I25369,g24891);
	nand 	XG14615 	(g27586,g26863,g24905,g24916,g24924);
	or 	XG14616 	(g29501,g27634,g28583);
	or 	XG14617 	(g29313,g27270,g28284);
	and 	XG14618 	(g29362,g28307,g27379);
	not 	XG14619 	(I25115,g25322);
	not 	XG14620 	(I25351,g24466);
	not 	XG14621 	(I25095,g25265);
	not 	XG14622 	(I25366,g24477);
	not 	XG14623 	(I25380,g24481);
	not 	XG14624 	(I25399,g24489);
	not 	XG14625 	(I25105,g25284);
	not 	XG14626 	(I25391,g24483);
	nor 	XG14627 	(g25776,g24369,g24380,g7166);
	nor 	XG14628 	(g25851,g24369,g24380,g4311);
	and 	XG14629 	(g30003,g9021,g28149);
	nand 	XG14630 	(g24792,I23951,I23950);
	and 	XG14631 	(g27146,g1648,g8187,g26148);
	or 	XG14632 	(g28068,g21838,g27310);
	or 	XG14633 	(g30369,g18439,g30066);
	and 	XG14634 	(g28214,g26625,g27731);
	and 	XG14635 	(g28234,g26686,g27877);
	and 	XG14636 	(g28136,g23135,g27382);
	or 	XG14637 	(g28098,g22016,g27683);
	and 	XG14638 	(g29637,g29134,g2533);
	or 	XG14639 	(g30366,g18417,g30122);
	and 	XG14640 	(g29940,g28758,g1740);
	or 	XG14641 	(g28104,g22108,g27697);
	nand 	XG14642 	(g27577,g25765,g24988,g25002,g25019);
	and 	XG14643 	(g29535,g28871,g2303);
	and 	XG14644 	(g28251,g23662,g27826);
	or 	XG14645 	(g28064,g21781,g27298);
	or 	XG14646 	(g28095,g21970,g27674);
	and 	XG14647 	(g27209,g2051,g8365,g26213);
	and 	XG14648 	(g29882,g29151,g2361);
	and 	XG14649 	(g29512,g28793,g2161);
	and 	XG14650 	(g27668,g25917,g1367);
	or 	XG14651 	(g27122,g25917,g22537);
	or 	XG14652 	(g30352,g18340,g30094);
	not 	XG14653 	(g28709,I27192);
	nand 	XG14654 	(g27593,g26861,g24906,g24950,g24972);
	and 	XG14655 	(g28213,g23380,g27720);
	or 	XG14656 	(g30378,g18487,g30125);
	and 	XG14657 	(g29577,g28946,g2441);
	and 	XG14658 	(g28133,g23108,g27367);
	and 	XG14659 	(g29870,g29130,g2421);
	and 	XG14660 	(g29854,g29092,g2197);
	and 	XG14661 	(g29585,g28920,g1756);
	and 	XG14662 	(g29587,g28935,g2181);
	and 	XG14663 	(g28217,g23391,g27733);
	or 	XG14664 	(g30364,g18411,g30086);
	and 	XG14665 	(g29838,g29044,g1636);
	or 	XG14666 	(g28091,g21913,g27665);
	and 	XG14667 	(g29688,g28713,g2509);
	and 	XG14668 	(g29683,g29046,g1821);
	or 	XG14669 	(g28103,g22097,g27696);
	and 	XG14670 	(g28312,g26608,g27828);
	and 	XG14671 	(g29943,g28765,g2165);
	and 	XG14672 	(g28148,g26093,g27355);
	and 	XG14673 	(g29662,g29049,g1848);
	and 	XG14674 	(g27040,g26226,g6573,g6565,g7812);
	or 	XG14675 	(g30300,g27252,g28246);
	or 	XG14676 	(g29486,g27595,g28537);
	or 	XG14677 	(g29496,g27615,g28567);
	or 	XG14678 	(g30314,g27266,g28268);
	or 	XG14679 	(g30307,g27260,g28256);
	or 	XG14680 	(g29489,g27601,g28550);
	nand 	XG14681 	(g25215,I24385,I24384);
	and 	XG14682 	(g28466,g17637,g27960);
	and 	XG14683 	(g28572,g15669,g27829);
	and 	XG14684 	(g29804,g29014,g1592);
	and 	XG14685 	(g29686,g29057,g2246);
	and 	XG14686 	(g29868,g29128,g2227);
	and 	XG14687 	(g29687,g29097,g2407);
	and 	XG14688 	(g29551,g28867,g2173);
	and 	XG14689 	(g29605,g28973,g2445);
	and 	XG14690 	(g28289,g26575,g27734);
	and 	XG14691 	(g29869,g29129,g2331);
	or 	XG14692 	(g28101,g22062,g27691);
	or 	XG14693 	(g30365,g18412,g30158);
	and 	XG14694 	(g27714,g26171,g26424,g25195,g22384);
	and 	XG14695 	(g27762,g26218,g26424,g25226,g22472);
	and 	XG14696 	(g29621,g28994,g2449);
	and 	XG14697 	(g28243,g23423,g27879);
	and 	XG14698 	(g29603,g29060,g2265);
	nand 	XG14699 	(g27468,g26852,g24925,g24932,g24951);
	and 	XG14700 	(g27727,g26195,g26424,g25211,g22432);
	and 	XG14701 	(g27817,g26236,g26424,g25245,g22498);
	and 	XG14702 	(g27162,g2208,g8259,g26171);
	and 	XG14703 	(g29553,g28911,g2437);
	and 	XG14704 	(g29895,g29170,g2495);
	or 	XG14705 	(g28100,g22051,g27690);
	not 	XG14706 	(g28147,I26654);
	and 	XG14707 	(g29619,g29060,g2269);
	and 	XG14708 	(g28557,g15647,g27772);
	and 	XG14709 	(g28494,g17741,g27973);
	or 	XG14710 	(g30371,g18445,g30099);
	and 	XG14711 	(g29664,g29060,g2273);
	and 	XG14712 	(g28112,g26162,g27352);
	or 	XG14713 	(g30304,g27259,g28255);
	or 	XG14714 	(g30311,g27265,g28265);
	and 	XG14715 	(g28218,g26645,g27768);
	and 	XG14716 	(g29615,g29049,g1844);
	and 	XG14717 	(g28200,g11383,g27652);
	and 	XG14718 	(g29665,g28696,g2375);
	not 	XG14719 	(g26718,g25168);
	and 	XG14720 	(g27210,g2476,g8373,g26218);
	or 	XG14721 	(g28094,g21959,g27673);
	and 	XG14722 	(g29840,g29056,g2153);
	and 	XG14723 	(g28229,g17213,g27345);
	or 	XG14724 	(g27261,g25996,g24544);
	and 	XG14725 	(g28495,g12465,g27012);
	and 	XG14726 	(g28111,g22716,g27343);
	or 	XG14727 	(g28065,g21792,g27299);
	and 	XG14728 	(g28242,g23626,g27769);
	and 	XG14729 	(g29600,g29049,g1840);
	and 	XG14730 	(g29851,g29079,g1668);
	not 	XG14731 	(I26409,g26187);
	not 	XG14732 	(I26406,g26187);
	and 	XG14733 	(g29710,g29094,g2380);
	or 	XG14734 	(g28062,g21746,g27288);
	or 	XG14735 	(g29238,g18292,g28178);
	and 	XG14736 	(g28130,g23063,g27353);
	and 	XG14737 	(g27658,g25786,g22491);
	and 	XG14738 	(g27039,g26223,g5535,g5527,g7738);
	or 	XG14739 	(g30372,g18446,g30110);
	or 	XG14740 	(g28067,g21827,g27309);
	and 	XG14741 	(g28467,g12295,g26993);
	or 	XG14742 	(g29482,g27588,g28524);
	or 	XG14743 	(g29488,g27600,g28547);
	and 	XG14744 	(g29582,g28608,g27766);
	not 	XG14745 	(g29961,g28892);
	not 	XG14746 	(g29920,g28824);
	and 	XG14747 	(g28205,g16746,g27516);
	and 	XG14748 	(g27073,g26281,g3881,g3873,g7121);
	or 	XG14749 	(g28097,g22005,g27682);
	or 	XG14750 	(g30363,g18407,g30121);
	nand 	XG14751 	(g25236,I24416,I24415);
	and 	XG14752 	(g29566,g28907,g2307);
	or 	XG14753 	(g29485,g27594,g28535);
	or 	XG14754 	(g29495,g27614,g28563);
	and 	XG14755 	(g29636,g29097,g2403);
	or 	XG14756 	(g27037,g26171,g26195,g26218,g26236);
	not 	XG14757 	(g27009,g25911);
	and 	XG14758 	(g28488,g17713,g27969);
	nand 	XG14759 	(g27796,g26171,g26424,g25263,g21228);
	nand 	XG14760 	(g27933,g26236,g26424,g25356,g21228);
	nand 	XG14761 	(g27903,g26218,g26424,g25316,g21228);
	nand 	XG14762 	(g27854,g26195,g26424,g25283,g21228);
	and 	XG14763 	(g29649,g28678,g2241);
	and 	XG14764 	(g29547,g28857,g1748);
	or 	XG14765 	(g30353,g18355,g30095);
	or 	XG14766 	(g30370,g18440,g30135);
	not 	XG14767 	(g30297,g28758);
	not 	XG14768 	(g29905,g28783);
	not 	XG14769 	(g29999,g28973);
	not 	XG14770 	(g29944,g28911);
	or 	XG14771 	(g30367,g18418,g30133);
	and 	XG14772 	(g28199,g16684,g27479);
	and 	XG14773 	(g29620,g29097,g2399);
	and 	XG14774 	(g29855,g29093,g2287);
	or 	XG14775 	(g28061,g21735,g27287);
	and 	XG14776 	(g28233,g23411,g27827);
	or 	XG14777 	(g30351,g18339,g30084);
	not 	XG14778 	(g29977,g28920);
	not 	XG14779 	(g29939,g28857);
	not 	XG14780 	(g30074,g29046);
	not 	XG14781 	(g29994,g29049);
	not 	XG14782 	(g30065,g29049);
	not 	XG14783 	(g30016,g29049);
	or 	XG14784 	(g28092,g21924,g27666);
	not 	XG14785 	(I26799,g27660);
	and 	XG14786 	(g27988,g23941,g26781);
	and 	XG14787 	(g29969,g20509,g28121);
	and 	XG14788 	(g30091,g20716,g28127);
	and 	XG14789 	(g29985,g20532,g28127);
	and 	XG14790 	(g30080,g20674,g28121);
	and 	XG14791 	(g27541,g23334,g26278);
	and 	XG14792 	(g27992,g23964,g26800);
	and 	XG14793 	(g29381,g19399,g28135);
	and 	XG14794 	(g29380,g19396,g28134);
	and 	XG14795 	(g29629,g19779,g28211);
	and 	XG14796 	(g29377,g19387,g28132);
	and 	XG14797 	(g29613,g19763,g28208);
	and 	XG14798 	(g27553,g23353,g26293);
	and 	XG14799 	(g31238,g20053,g29583);
	and 	XG14800 	(g25096,g20560,g23778);
	and 	XG14801 	(g29521,g28824,g1744);
	and 	XG14802 	(g29865,g29115,g1802);
	and 	XG14803 	(g29509,g28755,g1600);
	and 	XG14804 	(g29645,g29018,g1714);
	and 	XG14805 	(g28201,g16720,g27499);
	and 	XG14806 	(g28261,g23695,g27878);
	and 	XG14807 	(g29511,g28783,g1736);
	nand 	XG14808 	(g24798,I23963,I23962);
	and 	XG14809 	(g29538,g28914,g2563);
	or 	XG14810 	(g27108,g25911,g22522);
	and 	XG14811 	(g27664,g25911,g1024);
	and 	XG14812 	(g29731,g29118,g2089);
	or 	XG14813 	(g30333,g21699,g29834);
	and 	XG14814 	(g29853,g29081,g1862);
	and 	XG14815 	(g28143,g26083,g27344);
	and 	XG14816 	(g29573,g28892,g1752);
	and 	XG14817 	(g27217,g2610,g8418,g26236);
	and 	XG14818 	(g29584,g29018,g1706);
	or 	XG14819 	(g27248,g25953,g24880);
	or 	XG14820 	(g27241,g25984,g24584);
	and 	XG14821 	(g29926,g28736,g1604);
	and 	XG14822 	(g29964,g28830,g2008);
	and 	XG14823 	(g28226,g26667,g27825);
	nor 	XG14824 	(g31294,g29660,g11326);
	and 	XG14825 	(g29839,g29045,g1728);
	and 	XG14826 	(g29631,g28656,g1682);
	and 	XG14827 	(g27186,g2342,g8316,g26195);
	and 	XG14828 	(g29648,g29121,g2112);
	and 	XG14829 	(g28125,g26209,g27381);
	not 	XG14830 	(g29955,g28950);
	not 	XG14831 	(g30022,g29001);
	and 	XG14832 	(g30566,g29507,g26247);
	or 	XG14833 	(g30456,g21869,g29378);
	or 	XG14834 	(g31894,g21870,g30671);
	and 	XG14835 	(g29646,g28675,g1816);
	and 	XG14836 	(g29574,g28931,g2016);
	and 	XG14837 	(g27121,g26326,g136);
	and 	XG14838 	(g29852,g29080,g1772);
	and 	XG14839 	(g29601,g28955,g1890);
	not 	XG14840 	(g30102,g29157);
	not 	XG14841 	(g30055,g29157);
	not 	XG14842 	(g30068,g29157);
	not 	XG14843 	(g30113,g29154);
	not 	XG14844 	(g29983,g28977);
	not 	XG14845 	(g30040,g29025);
	and 	XG14846 	(g29514,g28780,g1608);
	or 	XG14847 	(g27244,g25995,g24652);
	not 	XG14848 	(g29995,g28955);
	not 	XG14849 	(g30303,g28786);
	and 	XG14850 	(g29602,g28962,g2020);
	not 	XG14851 	(g29976,g29018);
	not 	XG14852 	(g30052,g29018);
	not 	XG14853 	(g29993,g29018);
	not 	XG14854 	(g30063,g29015);
	not 	XG14855 	(g29925,g28820);
	not 	XG14856 	(g29960,g28885);
	not 	XG14857 	(g29996,g28962);
	not 	XG14858 	(g29941,g28900);
	and 	XG14859 	(g27765,g25886,g4146);
	not 	XG14860 	(g29929,g28914);
	not 	XG14861 	(g29312,g28877);
	and 	XG14862 	(g29563,g28853,g1616);
	not 	XG14863 	(g29927,g28861);
	not 	XG14864 	(g29978,g28927);
	and 	XG14865 	(g27822,g25893,g4157);
	not 	XG14866 	(g27320,I26004);
	and 	XG14867 	(g29617,g28987,g2024);
	and 	XG14868 	(g27686,g25849,g1291);
	not 	XG14869 	(g30053,g29121);
	not 	XG14870 	(g30037,g29121);
	not 	XG14871 	(g30087,g29121);
	not 	XG14872 	(g30097,g29118);
	not 	XG14873 	(g30018,g28987);
	not 	XG14874 	(g29963,g28931);
	not 	XG14875 	(g29893,g28755);
	not 	XG14876 	(g30292,g28736);
	and 	XG14877 	(g28585,g10530,g27063);
	not 	XG14878 	(g29911,g28780);
	not 	XG14879 	(g29948,g28853);
	and 	XG14880 	(g27678,g25830,g947);
	and 	XG14881 	(g29524,g28864,g2004);
	not 	XG14882 	(g29921,g28864);
	not 	XG14883 	(g30310,g28830);
	or 	XG14884 	(g29276,g18709,g28616);
	and 	XG14885 	(g29532,g28861,g1878);
	and 	XG14886 	(g29867,g29117,g1996);
	and 	XG14887 	(g29638,g29025,g2583);
	and 	XG14888 	(g29685,g28711,g2084);
	or 	XG14889 	(g30362,g18392,g30120);
	nand 	XG14890 	(g25199,I24365,I24364);
	and 	XG14891 	(g31271,g23300,g29706);
	or 	XG14892 	(g30349,g18333,g30051);
	and 	XG14893 	(g29599,g29018,g1710);
	or 	XG14894 	(g30377,g18472,g30124);
	or 	XG14895 	(g30387,g18524,g30151);
	and 	XG14896 	(g29661,g29015,g1687);
	and 	XG14897 	(g29709,g29121,g2116);
	and 	XG14898 	(g30670,g29359,g11330);
	or 	XG14899 	(g30360,g18386,g30145);
	or 	XG14900 	(g30361,g18391,g30109);
	and 	XG14901 	(g29684,g29085,g1982);
	and 	XG14902 	(g29530,g28820,g1612);
	or 	XG14903 	(g30348,g18329,g30083);
	and 	XG14904 	(g29633,g29085,g1978);
	and 	XG14905 	(g29951,g28786,g1874);
	or 	XG14906 	(g29279,g18741,g28442);
	and 	XG14907 	(g31527,g29343,g7553);
	and 	XG14908 	(g29568,g28950,g2571);
	and 	XG14909 	(g29634,g29121,g2108);
	or 	XG14910 	(g30356,g18365,g30096);
	and 	XG14911 	(g29667,g29157,g2671);
	or 	XG14912 	(g30355,g18360,g30131);
	or 	XG14913 	(g29233,g18234,g28171);
	or 	XG14914 	(g30376,g18471,g30112);
	or 	XG14915 	(g30368,g18435,g30098);
	and 	XG14916 	(g29894,g29169,g2070);
	or 	XG14917 	(g30354,g18359,g30064);
	and 	XG14918 	(g29517,g28827,g1870);
	and 	XG14919 	(g29586,g28927,g1886);
	and 	XG14920 	(g32053,g31509,g14176);
	nor 	XG14921 	(g32296,g12259,g31509,g9044);
	or 	XG14922 	(g30383,g18513,g30138);
	and 	XG14923 	(g29589,g28977,g2575);
	or 	XG14924 	(g30386,g18523,g30139);
	and 	XG14925 	(g29733,g29157,g2675);
	or 	XG14926 	(g30375,g18466,g30149);
	and 	XG14927 	(g29549,g28900,g2012);
	and 	XG14928 	(g29616,g29085,g1974);
	and 	XG14929 	(g29622,g29001,g2579);
	or 	XG14930 	(g30357,g18366,g30107);
	or 	XG14931 	(g30335,g18174,g29746);
	not 	XG14932 	(g32201,g31509);
	and 	XG14933 	(g31523,g29333,g7528);
	and 	XG14934 	(g29572,g28885,g1620);
	or 	XG14935 	(g31866,g18142,g31252);
	and 	XG14936 	(g27564,g23378,g26305);
	and 	XG14937 	(g29708,g29082,g1955);
	and 	XG14938 	(g29712,g28726,g2643);
	or 	XG14939 	(g30380,g18492,g30161);
	or 	XG14940 	(g30374,g18465,g30078);
	or 	XG14941 	(g30359,g18385,g30075);
	or 	XG14942 	(g30381,g18497,g30126);
	and 	XG14943 	(g29866,g29116,g1906);
	or 	XG14944 	(g27253,g26052,g24661);
	and 	XG14945 	(g31149,g23021,g29508);
	or 	XG14946 	(g31014,g28160,g29367);
	and 	XG14947 	(g29984,g28877,g2567);
	or 	XG14948 	(g30379,g18491,g30089);
	or 	XG14949 	(g31247,g13324,g29513);
	and 	XG14950 	(g27997,g23995,g26813);
	and 	XG14951 	(g29884,g29153,g2555);
	and 	XG14952 	(g29652,g29157,g2667);
	nand 	XG14953 	(g25271,I24463,I24462);
	and 	XG14954 	(g29740,g29154,g2648);
	and 	XG14955 	(g29881,g29150,g2040);
	and 	XG14956 	(g29880,g29149,g1936);
	or 	XG14957 	(g30350,g18334,g30118);
	or 	XG14958 	(g31221,g28204,g29494);
	or 	XG14959 	(g30384,g18517,g30101);
	nand 	XG14960 	(g24807,I23980,I23979);
	and 	XG14961 	(g29907,g29177,g2629);
	and 	XG14962 	(g27995,g23985,g26809);
	or 	XG14963 	(g30373,g18461,g30111);
	and 	XG14964 	(g29663,g28693,g1950);
	and 	XG14965 	(g32019,g22358,g30579);
	not 	XG14966 	(g31013,g29679);
	or 	XG14967 	(g29237,g18289,g28185);
	and 	XG14968 	(g29896,g29171,g2599);
	not 	XG14969 	(g30325,I28576);
	not 	XG14970 	(g31227,g29744);
	not 	XG14971 	(I28913,g30322);
	or 	XG14972 	(g27236,g25974,g24620);
	or 	XG14973 	(g30336,g18203,g29324);
	or 	XG14974 	(g29232,g18231,g28183);
	or 	XG14975 	(g27271,g26053,g24547);
	nand 	XG14976 	(g24760,I23919,I23918);
	or 	XG14977 	(g29278,g18740,g28626);
	or 	XG14978 	(g29277,g18710,g28440);
	nand 	XG14979 	(g25258,I24440,I24439);
	not 	XG14980 	(g31239,g29916);
	or 	XG14981 	(g31668,g28558,g29924);
	or 	XG14982 	(g29234,g18239,g28415);
	and 	XG14983 	(g27981,g23924,g26751);
	not 	XG14984 	(g29912,g28827);
	not 	XG14985 	(g29950,g28896);
	not 	XG14986 	(g30076,g29085);
	not 	XG14987 	(g30036,g29085);
	not 	XG14988 	(g30017,g29085);
	not 	XG14989 	(g30085,g29082);
	or 	XG14990 	(g29231,g18229,g28301);
	or 	XG14991 	(g30385,g18518,g30172);
	or 	XG14992 	(g30382,g18498,g30137);
	or 	XG14993 	(g30358,g18381,g30108);
	and 	XG14994 	(g30023,g20570,g28508);
	and 	XG14995 	(g29383,g19412,g28138);
	and 	XG14996 	(g29644,g19794,g28216);
	and 	XG14997 	(g29630,g19781,g28212);
	and 	XG14998 	(g30607,g18989,g30291);
	and 	XG14999 	(g30600,g18975,g30287);
	and 	XG15000 	(g32197,g20088,g31144);
	and 	XG15001 	(g29564,g28896,g1882);
	nand 	XG15002 	(g31262,g11679,g29916,g767);
	and 	XG15003 	(g30936,g29916,g8830);
	and 	XG15004 	(g30612,g29597,g26338);
	and 	XG15005 	(g30918,g29707,g8681);
	or 	XG15006 	(g29236,g18287,g28313);
	or 	XG15007 	(g29239,g18297,g28427);
	nor 	XG15008 	(g31134,g24732,g29679,g8033);
	and 	XG15009 	(g30577,g29679,g26267);
	or 	XG15010 	(g31020,g28164,g29375);
	or 	XG15011 	(g30342,g18261,g29330);
	or 	XG15012 	(g31964,g14544,g31654);
	not 	XG15013 	(g29897,I28128);
	and 	XG15014 	(g32040,g31243,g14122);
	or 	XG15015 	(g31670,g28573,g29937);
	or 	XG15016 	(g32155,g29475,g30935);
	and 	XG15017 	(g30731,g29361,g11374);
	and 	XG15018 	(g30730,g29778,g26346);
	nor 	XG15019 	(g31233,g24825,g29778,g8522);
	or 	XG15020 	(g31277,g28285,g29570);
	or 	XG15021 	(g31474,g13583,g29668);
	not 	XG15022 	(g31138,g29778);
	and 	XG15023 	(g31069,g14150,g29793);
	not 	XG15024 	(g31848,g29385);
	not 	XG15025 	(g31849,g29385);
	not 	XG15026 	(g31805,g29385);
	not 	XG15027 	(g31798,g29385);
	not 	XG15028 	(g31813,g29385);
	not 	XG15029 	(g31799,g29385);
	not 	XG15030 	(g31852,g29385);
	not 	XG15031 	(g31808,g29385);
	not 	XG15032 	(g31809,g29385);
	not 	XG15033 	(g31836,g29385);
	not 	XG15034 	(g31853,g29385);
	not 	XG15035 	(g31822,g29385);
	not 	XG15036 	(g31837,g29385);
	not 	XG15037 	(g31830,g29385);
	not 	XG15038 	(g31842,g29385);
	not 	XG15039 	(g31816,g29385);
	not 	XG15040 	(g31823,g29385);
	not 	XG15041 	(g31817,g29385);
	not 	XG15042 	(g31810,g29385);
	not 	XG15043 	(g31843,g29385);
	not 	XG15044 	(g31831,g29385);
	not 	XG15045 	(g31856,g29385);
	not 	XG15046 	(g31857,g29385);
	not 	XG15047 	(g31802,g29385);
	not 	XG15048 	(g31850,g29385);
	not 	XG15049 	(g31811,g29385);
	not 	XG15050 	(g31826,g29385);
	not 	XG15051 	(g31803,g29385);
	not 	XG15052 	(g31827,g29385);
	not 	XG15053 	(g31846,g29385);
	not 	XG15054 	(g31820,g29385);
	not 	XG15055 	(g31851,g29385);
	not 	XG15056 	(g31847,g29385);
	not 	XG15057 	(g31840,g29385);
	not 	XG15058 	(g31796,g29385);
	not 	XG15059 	(g31797,g29385);
	not 	XG15060 	(g31834,g29385);
	not 	XG15061 	(g31821,g29385);
	not 	XG15062 	(g31806,g29385);
	not 	XG15063 	(g31835,g29385);
	not 	XG15064 	(g31841,g29385);
	not 	XG15065 	(g31807,g29385);
	not 	XG15066 	(g31814,g29385);
	not 	XG15067 	(g31800,g29385);
	not 	XG15068 	(g31815,g29385);
	not 	XG15069 	(g31838,g29385);
	not 	XG15070 	(g31839,g29385);
	not 	XG15071 	(g31854,g29385);
	not 	XG15072 	(g31801,g29385);
	not 	XG15073 	(g31818,g29385);
	not 	XG15074 	(g31819,g29385);
	not 	XG15075 	(g31855,g29385);
	not 	XG15076 	(g31824,g29385);
	not 	XG15077 	(g31844,g29385);
	not 	XG15078 	(g31858,g29385);
	not 	XG15079 	(g31825,g29385);
	not 	XG15080 	(g31859,g29385);
	not 	XG15081 	(g31832,g29385);
	not 	XG15082 	(g31845,g29385);
	not 	XG15083 	(g31828,g29385);
	not 	XG15084 	(g31829,g29385);
	not 	XG15085 	(g31812,g29385);
	not 	XG15086 	(g31833,g29385);
	not 	XG15087 	(g31804,g29385);
	not 	XG15088 	(I27543,g28187);
	not 	XG15089 	(I28062,g29194);
	not 	XG15090 	(g29474,I27758);
	or 	XG15091 	(g27980,g26131,g26105);
	or 	XG15092 	(g27972,g26105,g26131);
	not 	XG15093 	(g26990,g26105);
	not 	XG15094 	(g27977,g26105);
	not 	XG15095 	(g26973,g26105);
	not 	XG15096 	(g27142,g26105);
	not 	XG15097 	(g27004,g26131);
	not 	XG15098 	(g26987,g26131);
	not 	XG15099 	(g27155,g26131);
	not 	XG15100 	(g27985,g26131);
	nand 	XG15101 	(g27282,g479,g26248,g26269,g11192);
	nor 	XG15102 	(g28340,g26339,g27439);
	and 	XG15103 	(I27508,g28033,g24083,g24082,g19935);
	and 	XG15104 	(I27513,g28034,g24090,g24089,g19984);
	not 	XG15105 	(g28326,g27414);
	and 	XG15106 	(g28035,I26531,I26530,g24103);
	and 	XG15107 	(I27539,g24137,g24136,g24135,g28040);
	and 	XG15108 	(I27534,g24130,g24129,g24128,g28039);
	and 	XG15109 	(I27519,g24109,g24108,g24107,g28036);
	and 	XG15110 	(I27524,g24116,g24115,g24114,g28037);
	and 	XG15111 	(I27529,g24123,g24122,g24121,g28038);
	not 	XG15112 	(g27402,I26100);
	nor 	XG15113 	(g28476,g26547,g27627);
	nor 	XG15114 	(g28521,g26604,g27649);
	nand 	XG15115 	(g27582,g26105,g26131,g10857);
	not 	XG15116 	(g26510,I25369);
	and 	XG15117 	(I27503,g28032,g24076,g24075,g19890);
	nor 	XG15118 	(g28491,g27617,g8114);
	nor 	XG15119 	(g28482,g27617,g3522);
	nand 	XG15120 	(g29186,g4507,g27051);
	and 	XG15121 	(g31142,g30039,g2527);
	and 	XG15122 	(g31147,g30054,g12286);
	or 	XG15123 	(g29479,g28116,g28113);
	nand 	XG15124 	(g28888,g8139,g27738);
	and 	XG15125 	(g28253,g27700,g23719);
	or 	XG15126 	(g28059,g18276,g27042);
	or 	XG15127 	(g30081,g11366,g28454);
	or 	XG15128 	(g31007,g28159,g29364);
	or 	XG15129 	(g29848,g26077,g28260);
	and 	XG15130 	(g31776,g29385,g21329);
	or 	XG15131 	(g29892,g26120,g28300);
	or 	XG15132 	(g29484,g22191,g28124);
	nor 	XG15133 	(g28981,g27999,g9234);
	nor 	XG15134 	(g28953,g27999,g5170);
	not 	XG15135 	(g26834,I25552);
	nor 	XG15136 	(g29193,g7812,g26994,g9529);
	nor 	XG15137 	(g28106,g26994,g7812);
	or 	XG15138 	(g31319,g28324,g29612);
	or 	XG15139 	(g31472,g28352,g29642);
	or 	XG15140 	(g29776,g22846,g28225);
	or 	XG15141 	(g31307,g28311,g29596);
	nand 	XG15142 	(g28990,g8310,g27882);
	or 	XG15143 	(g28186,g27146,g27161,g27185,g27209);
	and 	XG15144 	(g28290,g27759,g23780);
	and 	XG15145 	(g28637,g27011,g22399);
	or 	XG15146 	(g30163,g28523,g23381);
	nand 	XG15147 	(g28363,g13593,g27064);
	nand 	XG15148 	(g28376,g13620,g27064);
	nand 	XG15149 	(g28406,g13675,g27064);
	nand 	XG15150 	(g28391,g13637,g27064);
	nand 	XG15151 	(g28395,g13655,g27074);
	nand 	XG15152 	(g28381,g13621,g27074);
	nand 	XG15153 	(g28410,g13679,g27074);
	nand 	XG15154 	(g28421,g13715,g27074);
	or 	XG15155 	(g29480,g22172,g28115);
	nor 	XG15156 	(g29167,g26994,g9576);
	nor 	XG15157 	(g29146,g26994,g6565);
	or 	XG15158 	(g29792,g28244,g28235);
	or 	XG15159 	(g30176,g28531,g23392);
	not 	XG15160 	(g27961,g26816);
	and 	XG15161 	(g31210,g30100,g2509);
	or 	XG15162 	(g29849,g28273,g26049);
	nor 	XG15163 	(g29173,g7704,g27999,g9259);
	nor 	XG15164 	(g29187,g27999,g7704);
	nor 	XG15165 	(g29370,g28599,g28585);
	not 	XG15166 	(g26825,I25541);
	nand 	XG15167 	(g28965,g8255,g27882);
	nand 	XG15168 	(g28934,g14641,g27882);
	nor 	XG15169 	(g29184,g26994,g9631);
	nor 	XG15170 	(g29181,g26994,g6573);
	nand 	XG15171 	(g28856,g8093,g27738);
	nand 	XG15172 	(g28823,g14565,g27738);
	not 	XG15173 	(g26859,I25591);
	or 	XG15174 	(g30141,g16844,g28499);
	not 	XG15175 	(g26850,I25576);
	nand 	XG15176 	(g28923,g8195,g27775);
	and 	XG15177 	(g28263,g27711,g23747);
	not 	XG15178 	(g27929,I26448);
	and 	XG15179 	(g31169,g30079,g10083);
	not 	XG15180 	(g26835,I25555);
	and 	XG15181 	(g31790,g29385,g21299);
	or 	XG15182 	(g31375,g28339,g29628);
	not 	XG15183 	(I26195,g26260);
	nor 	XG15184 	(g28031,I26523,I26522,g21209);
	or 	XG15185 	(g28057,g18218,g27033);
	or 	XG15186 	(g29692,g10873,g28197);
	not 	XG15187 	(g28559,g27700);
	not 	XG15188 	(g28590,g27724);
	nor 	XG15189 	(g29007,g28010,g9269);
	nor 	XG15190 	(g28986,g28010,g5517);
	not 	XG15191 	(g25903,I25005);
	nor 	XG15192 	(g29107,g26977,g7791,g6203);
	nor 	XG15193 	(g29180,g26977,g9569);
	nor 	XG15194 	(g29175,g26977,g6227);
	nor 	XG15195 	(g29069,g28010,g9381);
	nor 	XG15196 	(g29034,g28010,g5527);
	not 	XG15197 	(g28575,g27711);
	not 	XG15198 	(g28604,g27759);
	not 	XG15199 	(g27881,I26430);
	not 	XG15200 	(I26516,g26824);
	or 	XG15201 	(g30115,g11449,g28489);
	not 	XG15202 	(I27677,g28156);
	and 	XG15203 	(g31152,g30067,g10039);
	or 	XG15204 	(g29502,g25871,g28139);
	and 	XG15205 	(g31788,g29385,g21352);
	not 	XG15206 	(g26817,g25242);
	or 	XG15207 	(g29864,g26086,g28272);
	nor 	XG15208 	(g28457,g27602,g7980);
	nor 	XG15209 	(g28452,g27602,g3161);
	and 	XG15210 	(g31186,g30088,g2375);
	nor 	XG15211 	(g28492,g27635,g7121,g3857);
	nor 	XG15212 	(g28483,g27635,g8080);
	nor 	XG15213 	(g28475,g27635,g3863);
	or 	XG15214 	(g28209,g27141,g27223);
	not 	XG15215 	(g28443,I26936);
	or 	XG15216 	(g29786,g28240,g22843);
	nor 	XG15217 	(g29070,g28020,g7766,g5857);
	or 	XG15218 	(g29756,g28223,g22717);
	nor 	XG15219 	(g29035,g28020,g9321);
	nor 	XG15220 	(g29012,g28020,g5863);
	nand 	XG15221 	(g28930,g8201,g27833);
	or 	XG15222 	(g29775,g28232,g25966);
	or 	XG15223 	(g30189,g28543,g23401);
	not 	XG15224 	(g26843,I25567);
	nor 	XG15225 	(g29072,g26977,g9402);
	nor 	XG15226 	(g29040,g26977,g6209);
	nor 	XG15227 	(g28414,g26347,g27467);
	and 	XG15228 	(g27395,g9077,g9187,g26314,g8046);
	and 	XG15229 	(g27421,g9077,g9187,g26314,g8038);
	and 	XG15230 	(g27416,g504,g9187,g26314,g8046);
	and 	XG15231 	(g27445,g504,g9187,g26314,g8038);
	or 	XG15232 	(g31001,g28151,g29360);
	nor 	XG15233 	(g29141,g27999,g9374);
	nor 	XG15234 	(g29104,g27999,g5188);
	and 	XG15235 	(g27474,g504,g518,g26314,g8038);
	and 	XG15236 	(g27494,g9077,g518,g26314,g8038);
	and 	XG15237 	(g27440,g504,g518,g26314,g8046);
	and 	XG15238 	(g27469,g9077,g518,g26314,g8046);
	nor 	XG15239 	(g28520,g27635,g8229);
	nor 	XG15240 	(g28515,g27635,g3881);
	nor 	XG15241 	(g29109,g26994,g9472);
	nor 	XG15242 	(g29077,g26994,g6555);
	not 	XG15243 	(I26508,g26814);
	nor 	XG15244 	(g29164,g28010,g9444);
	or 	XG15245 	(I26644,g27032,g27039,g27044,g27057);
	nor 	XG15246 	(g29142,g28010,g5535);
	and 	XG15247 	(g31131,g30020,g2393);
	and 	XG15248 	(g31141,g30038,g12224);
	or 	XG15249 	(g30103,g16731,g28477);
	nand 	XG15250 	(g28895,g8146,g27775);
	nand 	XG15251 	(g28860,g14586,g27775);
	not 	XG15252 	(I26581,g26942);
	nor 	XG15253 	(g28480,g27602,g8059);
	nor 	XG15254 	(g28469,g27602,g3171);
	nor 	XG15255 	(g29174,g28020,g9511);
	nor 	XG15256 	(g29165,g28020,g5881);
	or 	XG15257 	(g29735,g10898,g28202);
	and 	XG15258 	(g31778,g29385,g21369);
	not 	XG15259 	(I29207,g30293);
	not 	XG15260 	(I26503,g26811);
	not 	XG15261 	(g25771,I24920);
	and 	XG15262 	(g30564,g29385,g21358);
	nor 	XG15263 	(g28584,g27635,g7121);
	nor 	XG15264 	(g28540,g7121,g27635,g8125);
	nor 	XG15265 	(g28498,g27635,g8172);
	or 	XG15266 	(I26643,g27040,g27045,g27058,g27073);
	nor 	XG15267 	(g28493,g27635,g3873);
	not 	XG15268 	(g26648,g25115);
	not 	XG15269 	(I29211,g30298);
	and 	XG15270 	(g27669,g13278,g26840);
	not 	XG15271 	(I26584,g26943);
	or 	XG15272 	(g30104,g11427,g28478);
	or 	XG15273 	(g29148,g26606,g27651);
	and 	XG15274 	(g31759,g29385,g21291);
	nor 	XG15275 	(g29145,g26994,g7812,g6549);
	nor 	XG15276 	(g29005,g27999,g7704,g5164);
	nor 	XG15277 	(g29198,g28020,g7766);
	nor 	XG15278 	(g29183,g7766,g28020,g9392);
	nor 	XG15279 	(g29106,g28020,g9451);
	nor 	XG15280 	(g29071,g28020,g5873);
	nor 	XG15281 	(g28425,g26351,g27493);
	not 	XG15282 	(g26851,I25579);
	nand 	XG15283 	(g27273,g26105,g26131,g10504);
	and 	XG15284 	(g31787,g29385,g21281);
	and 	XG15285 	(g31777,g29385,g21343);
	not 	XG15286 	(g25220,I24396);
	not 	XG15287 	(g26862,I25598);
	not 	XG15288 	(g26870,I25606);
	not 	XG15289 	(I25511,g25073);
	not 	XG15290 	(I25514,g25073);
	not 	XG15291 	(g28380,g27064);
	not 	XG15292 	(g28241,g27064);
	nand 	XG15293 	(g28109,g25783,g27051);
	nand 	XG15294 	(g28131,g25838,g27051);
	and 	XG15295 	(g28114,g27051,g25869);
	not 	XG15296 	(I27401,g27051);
	not 	XG15297 	(g28250,g27074);
	not 	XG15298 	(g28399,g27074);
	not 	XG15299 	(I26578,g26941);
	not 	XG15300 	(I28185,g28803);
	not 	XG15301 	(I28199,g28803);
	not 	XG15302 	(I27927,g28803);
	not 	XG15303 	(I28174,g28803);
	not 	XG15304 	(I27941,g28803);
	not 	XG15305 	(I27954,g28803);
	not 	XG15306 	(I27970,g28803);
	not 	XG15307 	(I28162,g28803);
	and 	XG15308 	(g28158,g27037,g22763,g26424);
	not 	XG15309 	(g28274,I26799);
	and 	XG15310 	(g28153,g27031,g22763,g26424);
	or 	XG15311 	(g31293,g28299,g29582);
	or 	XG15312 	(g29716,g15856,g28199);
	nor 	XG15313 	(g29108,g26977,g6219);
	nor 	XG15314 	(g29144,g26977,g9518);
	nor 	XG15315 	(g28462,g27617,g3512);
	nor 	XG15316 	(g28470,g27617,g8021);
	nor 	XG15317 	(g28468,g27602,g10295,g3155);
	or 	XG15318 	(g29717,g10883,g28200);
	or 	XG15319 	(g29791,g22859,g28233);
	or 	XG15320 	(g30201,g28557,g23412);
	nor 	XG15321 	(g28519,g10295,g27602,g8011);
	nor 	XG15322 	(g28552,g27602,g10295);
	nor 	XG15323 	(g29006,g27999,g5180);
	nor 	XG15324 	(g29032,g27999,g9300);
	and 	XG15325 	(g28624,g27009,g22357);
	or 	XG15326 	(g29777,g28234,g28227);
	nor 	XG15327 	(g29189,g7791,g26977,g9462);
	nor 	XG15328 	(g29200,g26977,g7791);
	and 	XG15329 	(g25968,g20739,g25215);
	nor 	XG15330 	(g28481,g27617,g10323,g3506);
	or 	XG15331 	(g30127,g16805,g28494);
	and 	XG15332 	(g25787,g20887,g24792);
	or 	XG15333 	(g29487,g28133,g25815);
	and 	XG15334 	(g28280,g27724,g23761);
	nand 	XG15335 	(g28899,g14612,g27833);
	nand 	XG15336 	(g28958,g8249,g27833);
	or 	XG15337 	(g29476,g28112,g28108);
	and 	XG15338 	(g28302,g27817,g23809);
	nand 	XG15339 	(g29028,g8381,g27933);
	or 	XG15340 	(g30093,g11397,g28467);
	nor 	XG15341 	(g28510,g27617,g3530);
	nor 	XG15342 	(g28514,g27617,g8165);
	or 	XG15343 	(g29768,g28229,g22760);
	or 	XG15344 	(g30128,g11497,g28495);
	and 	XG15345 	(g31130,g30019,g12191);
	and 	XG15346 	(g31124,g29997,g2259);
	nor 	XG15347 	(g29033,g28010,g7738,g5511);
	nor 	XG15348 	(g28529,g10323,g27617,g8070);
	nor 	XG15349 	(g28568,g27617,g10323);
	or 	XG15350 	(g29879,g26096,g28289);
	nor 	XG15351 	(g28496,g27602,g3179);
	nor 	XG15352 	(g28509,g27602,g8107);
	nor 	XG15353 	(g29191,g28010,g7738);
	nor 	XG15354 	(g29179,g7738,g28010,g9311);
	and 	XG15355 	(g28282,g27727,g23762);
	or 	XG15356 	(g28191,g27162,g27186,g27210,g27217);
	nand 	XG15357 	(g28969,g8267,g27854);
	or 	XG15358 	(g28194,g27122,g22540);
	and 	XG15359 	(g28673,g27122,g1373);
	or 	XG15360 	(g29506,g25880,g28148);
	and 	XG15361 	(g31168,g30077,g2241);
	or 	XG15362 	(g29753,g22720,g28213);
	or 	XG15363 	(g30114,g16761,g28488);
	or 	XG15364 	(g30092,g16699,g28466);
	nand 	XG15365 	(I29261,g12046,g29485);
	nand 	XG15366 	(I29277,g12081,g29488);
	or 	XG15367 	(g29741,g15883,g28205);
	or 	XG15368 	(g29748,g28214,g28210);
	or 	XG15369 	(g29790,g28242,g25975);
	or 	XG15370 	(g29483,g28130,g25801);
	or 	XG15371 	(g29168,g26613,g27658);
	or 	XG15372 	(g29478,g22160,g28111);
	or 	XG15373 	(g29754,g28218,g28215);
	not 	XG15374 	(g27832,I26409);
	or 	XG15375 	(g29763,g22762,g28217);
	or 	XG15376 	(g31002,g28154,g29362);
	and 	XG15377 	(g31187,g30090,g10118);
	nand 	XG15378 	(I29269,g12050,g29486);
	and 	XG15379 	(g28292,g27762,g23781);
	not 	XG15380 	(g27737,g26718);
	nand 	XG15381 	(I29284,g12085,g29489);
	nand 	XG15382 	(I29313,g12154,g29501);
	not 	XG15383 	(I29225,g30311);
	not 	XG15384 	(I29218,g30304);
	not 	XG15385 	(I28548,g28147);
	or 	XG15386 	(g29802,g22871,g28243);
	and 	XG15387 	(g28266,g27714,g23748);
	not 	XG15388 	(g28615,g27817);
	not 	XG15389 	(g28593,g27727);
	or 	XG15390 	(g30214,g28572,g23424);
	or 	XG15391 	(g29904,g26146,g28312);
	not 	XG15392 	(g28606,g27762);
	not 	XG15393 	(g28579,g27714);
	or 	XG15394 	(g29801,g28251,g25987);
	not 	XG15395 	(I29221,g30307);
	not 	XG15396 	(I29228,g30314);
	not 	XG15397 	(I29214,g30300);
	or 	XG15398 	(g29490,g28136,g25832);
	not 	XG15399 	(I28241,g28709);
	not 	XG15400 	(g28126,g27122);
	not 	XG15401 	(I25869,g25851);
	not 	XG15402 	(I25882,g25776);
	not 	XG15403 	(g26549,I25391);
	not 	XG15404 	(g26026,I25105);
	not 	XG15405 	(g26576,I25399);
	not 	XG15406 	(g26519,I25380);
	not 	XG15407 	(g26488,I25366);
	not 	XG15408 	(g25997,I25095);
	not 	XG15409 	(g26400,I25351);
	not 	XG15410 	(g26055,I25115);
	not 	XG15411 	(I29242,g29313);
	or 	XG15412 	(g28096,g21997,g27988);
	nand 	XG15413 	(I29295,g12117,g29495);
	and 	XG15414 	(g31209,g30097,g2084);
	and 	XG15415 	(g31148,g30055,g2661);
	and 	XG15416 	(g31153,g30068,g12336);
	or 	XG15417 	(g28066,g21819,g27553);
	nand 	XG15418 	(g28976,g8273,g27903);
	and 	XG15419 	(g31185,g30087,g10114);
	and 	XG15420 	(g31123,g29994,g1834);
	and 	XG15421 	(g31128,g30016,g12187);
	or 	XG15422 	(g30340,g18245,g29377);
	or 	XG15423 	(g30346,g18303,g29381);
	nand 	XG15424 	(I29302,g12121,g29496);
	or 	XG15425 	(g30392,g18558,g30091);
	and 	XG15426 	(g31151,g30065,g10037);
	nand 	XG15427 	(g28906,g8150,g27796);
	nand 	XG15428 	(g28870,g14588,g27796);
	or 	XG15429 	(g30341,g18246,g29380);
	and 	XG15430 	(g31211,g30102,g10156);
	nand 	XG15431 	(g28938,g8205,g27796);
	or 	XG15432 	(g30389,g18554,g29969);
	and 	XG15433 	(g31222,g30113,g2643);
	nand 	XG15434 	(g28949,g14643,g27903);
	nand 	XG15435 	(g28997,g8324,g27903);
	not 	XG15436 	(I27235,g27320);
	not 	XG15437 	(I27238,g27320);
	or 	XG15438 	(g29734,g15872,g28201);
	or 	XG15439 	(g28063,g21773,g27541);
	or 	XG15440 	(g29813,g28261,g26020);
	and 	XG15441 	(g25977,g20875,g25236);
	or 	XG15442 	(g30338,g18240,g29613);
	nand 	XG15443 	(I29253,g12017,g29482);
	nand 	XG15444 	(g29004,g8330,g27933);
	or 	XG15445 	(g29504,g25875,g28143);
	or 	XG15446 	(g30390,g18555,g29985);
	nand 	XG15447 	(g28980,g14680,g27933);
	and 	XG15448 	(g31166,g30074,g1816);
	nand 	XG15449 	(g28945,g8211,g27854);
	nand 	XG15450 	(g28910,g14614,g27854);
	or 	XG15451 	(g29481,g28125,g28117);
	and 	XG15452 	(g28654,g27108,g1030);
	or 	XG15453 	(g28188,g27108,g22535);
	or 	XG15454 	(g29764,g28226,g28219);
	nor 	XG15455 	(g32424,g31294,g8721);
	or 	XG15456 	(g30339,g18244,g29629);
	or 	XG15457 	(g28099,g22043,g27992);
	or 	XG15458 	(g31867,g18175,g31238);
	and 	XG15459 	(g25803,g21024,g24798);
	or 	XG15460 	(g25616,g18172,g25096);
	not 	XG15461 	(g28120,g27108);
	or 	XG15462 	(g30391,g18557,g30080);
	and 	XG15463 	(g31948,g18884,g30670);
	and 	XG15464 	(g32425,g21604,g31668);
	and 	XG15465 	(g32169,g23046,g31014);
	and 	XG15466 	(g32207,g23323,g31221);
	and 	XG15467 	(g32254,g20379,g31247);
	and 	XG15468 	(g31145,g30052,g9970);
	and 	XG15469 	(g31139,g30036,g12221);
	and 	XG15470 	(g31129,g30017,g1968);
	and 	XG15471 	(g32034,g31239,g14124);
	nand 	XG15472 	(g33299,g12323,g32296,g608);
	and 	XG15473 	(g33124,g32296,g8945);
	and 	XG15474 	(g25817,g21163,g24807);
	or 	XG15475 	(g28093,g21951,g27981);
	or 	XG15476 	(g28069,g21865,g27564);
	and 	XG15477 	(g31150,g30063,g1682);
	and 	XG15478 	(g31962,g31013,g8033);
	or 	XG15479 	(g33035,g21872,g32019);
	not 	XG15480 	(g30931,I28913);
	not 	XG15481 	(I29371,g30325);
	or 	XG15482 	(g32037,g29329,g30566);
	and 	XG15483 	(g31122,g29993,g12144);
	and 	XG15484 	(g31120,g29976,g1700);
	or 	XG15485 	(g28102,g22089,g27995);
	or 	XG15486 	(g28105,g22135,g27997);
	or 	XG15487 	(g31865,g21709,g31149);
	and 	XG15488 	(g25961,g20682,g25199);
	or 	XG15489 	(g32395,g30049,g31523);
	and 	XG15490 	(g31146,g30053,g12285);
	and 	XG15491 	(g31140,g30037,g2102);
	not 	XG15492 	(g33258,g32296);
	or 	XG15493 	(g31864,g21703,g31271);
	or 	XG15494 	(g30388,g18534,g30023);
	or 	XG15495 	(g32978,g18145,g32197);
	or 	XG15496 	(g30347,g18304,g29383);
	and 	XG15497 	(g31167,g30076,g10080);
	or 	XG15498 	(g30345,g18302,g29644);
	or 	XG15499 	(g32399,g30062,g31527);
	or 	XG15500 	(g30344,g18298,g29630);
	and 	XG15501 	(g33126,g32201,g9044);
	or 	XG15502 	(g31870,g18262,g30607);
	and 	XG15503 	(g26022,g20751,g25271);
	or 	XG15504 	(g33235,g30982,g32040);
	and 	XG15505 	(g25814,g13323,g24760);
	and 	XG15506 	(g25989,g21012,g25258);
	and 	XG15507 	(g32011,g31134,g8287);
	and 	XG15508 	(g32173,g31134,g160);
	and 	XG15509 	(g31184,g30085,g1950);
	and 	XG15510 	(g33113,g22339,g31964);
	not 	XG15511 	(g32137,g31134);
	or 	XG15512 	(g31868,g18204,g30600);
	or 	XG15513 	(g32125,g29376,g30918);
	not 	XG15514 	(g32192,g31262);
	and 	XG15515 	(g31524,g20593,g29897);
	and 	XG15516 	(g32339,g20672,g31474);
	and 	XG15517 	(g31934,g18827,g31670);
	and 	XG15518 	(g31963,g18895,g30731);
	and 	XG15519 	(g33252,g20064,g32155);
	and 	XG15520 	(g32181,g19912,g31020);
	and 	XG15521 	(g32041,g31262,g13913);
	nor 	XG15522 	(g32212,g11083,g31262,g8859);
	or 	XG15523 	(g32094,g29363,g30612);
	and 	XG15524 	(g32190,g31233,g142);
	and 	XG15525 	(g32012,g31233,g8297);
	and 	XG15526 	(g32154,g14184,g31277);
	not 	XG15527 	(g32138,g31233);
	and 	XG15528 	(g32016,g31138,g8522);
	or 	XG15529 	(g32202,g13410,g31069);
	nand 	XG15530 	(g28512,g27142,g27155,g10857);
	nand 	XG15531 	(g28522,g27142,g26131,g10857);
	nand 	XG15532 	(g28516,g27155,g26105,g10857);
	and 	XG15533 	(g29208,I27539,I27538,g24138);
	and 	XG15534 	(g29203,I27514,I27513,g24095);
	and 	XG15535 	(g29202,I27509,I27508,g24088);
	and 	XG15536 	(g28652,g10288,g27282);
	nand 	XG15537 	(g28288,g27004,g26105,g10533);
	nand 	XG15538 	(g28271,g26990,g27004,g10533);
	nand 	XG15539 	(g28298,g26990,g26131,g10533);
	nand 	XG15540 	(g28259,g26973,g26987,g10504);
	nand 	XG15541 	(g28287,g26973,g26131,g10504);
	nand 	XG15542 	(g28270,g26987,g26105,g10504);
	nand 	XG15543 	(g28203,g27977,g27985,g12546);
	nand 	XG15544 	(g28206,g27985,g26105,g12546);
	nand 	XG15545 	(g28207,g27977,g26131,g12546);
	not 	XG15546 	(I26952,g27972);
	not 	XG15547 	(I26929,g27980);
	not 	XG15548 	(I28579,g29474);
	not 	XG15549 	(g29814,I28062);
	not 	XG15550 	(g29209,I27543);
	and 	XG15551 	(g32341,g23610,g31472);
	and 	XG15552 	(g31494,g23435,g29792);
	and 	XG15553 	(g31769,g23986,g30141);
	and 	XG15554 	(g31517,g23482,g29849);
	and 	XG15555 	(g29338,g22181,g29145);
	and 	XG15556 	(g31784,g24003,g30176);
	and 	XG15557 	(g31519,g23490,g29864);
	and 	XG15558 	(g32316,g23522,g31307);
	and 	XG15559 	(g31750,g23925,g30103);
	and 	XG15560 	(g31125,g22973,g29502);
	and 	XG15561 	(g31475,g23406,g29756);
	and 	XG15562 	(g32160,g22995,g31001);
	and 	XG15563 	(g31270,g23282,g29692);
	and 	XG15564 	(g32327,g23544,g31319);
	and 	XG15565 	(g31485,g23421,g29776);
	and 	XG15566 	(g31786,g24010,g30189);
	and 	XG15567 	(g31752,g23928,g30104);
	and 	XG15568 	(g29327,g22156,g29070);
	and 	XG15569 	(g31707,g23886,g30081);
	and 	XG15570 	(g31484,g23418,g29775);
	and 	XG15571 	(g31516,g23476,g29848);
	and 	XG15572 	(g31780,g23999,g30163);
	and 	XG15573 	(g29314,g22144,g29005);
	and 	XG15574 	(g29369,g22341,g28209);
	and 	XG15575 	(g29334,g18908,g29148);
	and 	XG15576 	(g31018,g22855,g29480);
	and 	XG15577 	(g31017,g22841,g29479);
	and 	XG15578 	(g29332,g22170,g29107);
	and 	XG15579 	(g31525,g23526,g29892);
	and 	XG15580 	(g32334,g23568,g31375);
	and 	XG15581 	(g31758,g23945,g30115);
	and 	XG15582 	(g32166,g23029,g31007);
	and 	XG15583 	(g31292,g23338,g29735);
	and 	XG15584 	(g31067,g22868,g29484);
	and 	XG15585 	(g31490,g23429,g29786);
	and 	XG15586 	(g30025,g23502,g28492);
	not 	XG15587 	(g29930,I28162);
	not 	XG15588 	(g29713,I27970);
	not 	XG15589 	(g29689,I27954);
	not 	XG15590 	(g29669,I27941);
	not 	XG15591 	(g29945,I28174);
	not 	XG15592 	(g29653,I27927);
	not 	XG15593 	(g29970,I28199);
	not 	XG15594 	(g29956,I28185);
	nor 	XG15595 	(g29503,g28250,g22763);
	nor 	XG15596 	(g29497,g28241,g22763);
	not 	XG15597 	(g28079,I26578);
	not 	XG15598 	(g29067,I27401);
	not 	XG15599 	(I28434,g28114);
	and 	XG15600 	(g30026,g25064,g28476);
	and 	XG15601 	(g30004,g25837,g28521);
	and 	XG15602 	(g29835,g24866,g28326);
	and 	XG15603 	(g29803,g26836,g28414);
	and 	XG15604 	(g29850,g24893,g28340);
	and 	XG15605 	(g29836,g26841,g28425);
	and 	XG15606 	(g28264,g27416,g1802,g7315);
	and 	XG15607 	(g29571,g11762,g28452);
	and 	XG15608 	(g29579,g7964,g28457);
	and 	XG15609 	(g29592,g11832,g28469);
	and 	XG15610 	(g29606,g8011,g28480);
	not 	XG15611 	(g26802,I25514);
	and 	XG15612 	(g30069,g12708,g29175);
	and 	XG15613 	(g30058,g12950,g29180);
	and 	XG15614 	(g31504,g10553,g29370);
	not 	XG15615 	(I26466,g26870);
	not 	XG15616 	(I26451,g26862);
	not 	XG15617 	(g26810,g25220);
	and 	XG15618 	(g28970,g27445,g26424,g25196,g17405);
	and 	XG15619 	(g28939,g27421,g26424,g25184,g17321);
	and 	XG15620 	(g29548,g28575,g1798);
	or 	XG15621 	(g32219,g29620,g31131);
	and 	XG15622 	(g29354,g28421,g4961);
	and 	XG15623 	(g29975,g10420,g28986);
	and 	XG15624 	(g29990,g9239,g29007);
	and 	XG15625 	(g29609,g11861,g28482);
	and 	XG15626 	(g29624,g8070,g28491);
	and 	XG15627 	(g29345,g28376,g4749);
	and 	XG15628 	(g30009,g10518,g29034);
	and 	XG15629 	(g30028,g9311,g29069);
	and 	XG15630 	(g28991,g27469,g26424,g25209,g14438);
	and 	XG15631 	(g28959,g27440,g26424,g25194,g17401);
	or 	XG15632 	(g30286,g28186,g28191);
	and 	XG15633 	(g29531,g28559,g1664);
	not 	XG15634 	(I26381,g26851);
	and 	XG15635 	(g29029,g27494,g26424,g25227,g14506);
	and 	XG15636 	(g28998,g27474,g26424,g25212,g17424);
	and 	XG15637 	(g30056,g12659,g29165);
	and 	XG15638 	(g30044,g12944,g29174);
	and 	XG15639 	(g29959,g12823,g28953);
	and 	XG15640 	(g29973,g9206,g28981);
	and 	XG15641 	(g30034,g10541,g29077);
	and 	XG15642 	(g30047,g9407,g29109);
	nand 	XG15643 	(g29719,g13739,g28406);
	nand 	XG15644 	(g29657,g13634,g28363);
	not 	XG15645 	(g28081,I26584);
	or 	XG15646 	(g32275,g29732,g31210);
	or 	XG15647 	(g32222,g29636,g31141);
	not 	XG15648 	(g31609,I29211);
	not 	XG15649 	(g27698,g26648);
	or 	XG15650 	(g28140,I26644,I26643);
	and 	XG15651 	(g29656,g11666,g28515);
	and 	XG15652 	(g29641,g14237,g28520);
	or 	XG15653 	(g32228,g29651,g31147);
	not 	XG15654 	(I26479,g25771);
	not 	XG15655 	(g27993,I26503);
	and 	XG15656 	(g28303,g27494,g2629,g7462);
	not 	XG15657 	(g31601,I29207);
	not 	XG15658 	(g28080,I26581);
	and 	XG15659 	(g29352,g28410,g4950);
	not 	XG15660 	(g27996,I26508);
	and 	XG15661 	(g30059,g12467,g28106);
	and 	XG15662 	(g30048,g12945,g29193);
	or 	XG15663 	(g28172,g27395,g27416,g27440,g27469);
	or 	XG15664 	(g28179,g27421,g27445,g27474,g27494);
	or 	XG15665 	(g32262,g29710,g31186);
	and 	XG15666 	(g29349,g28391,g4760);
	not 	XG15667 	(I26356,g26843);
	or 	XG15668 	(I26741,g27402,g22928,g22905,g22881);
	and 	XG15669 	(g28453,g10233,g27582);
	and 	XG15670 	(g29336,g28363,g4704);
	not 	XG15671 	(I28458,g28443);
	and 	XG15672 	(g29346,g28381,g4894);
	not 	XG15673 	(I26512,g26817);
	or 	XG15674 	(g32236,g29664,g31152);
	and 	XG15675 	(g29351,g28406,g4771);
	not 	XG15676 	(g29317,I27677);
	nand 	XG15677 	(g29737,g13779,g28421);
	nand 	XG15678 	(g29676,g13676,g28381);
	nand 	XG15679 	(g29694,g13709,g28391);
	nand 	XG15680 	(g29672,g13672,g28376);
	not 	XG15681 	(g28009,I26516);
	not 	XG15682 	(I27368,g27881);
	nand 	XG15683 	(g29722,g13742,g28410);
	nand 	XG15684 	(g29702,g13712,g28395);
	and 	XG15685 	(g29534,g22457,g28965);
	and 	XG15686 	(g29550,g22457,g28990);
	and 	XG15687 	(g29647,g22457,g28934);
	and 	XG15688 	(g29522,g22369,g28923);
	not 	XG15689 	(I25743,g25903);
	and 	XG15690 	(g29598,g22342,g28823);
	and 	XG15691 	(g29510,g22342,g28856);
	and 	XG15692 	(g29515,g22342,g28888);
	and 	XG15693 	(g29206,I27529,I27528,g24124);
	and 	XG15694 	(g29201,I27504,I27503,g24081);
	and 	XG15695 	(g29205,I27524,I27523,g24117);
	and 	XG15696 	(g29204,I27519,I27518,g24110);
	and 	XG15697 	(g29207,I27534,I27533,g24131);
	not 	XG15698 	(g27527,I26195);
	not 	XG15699 	(I26337,g26835);
	or 	XG15700 	(g32249,g29687,g31169);
	not 	XG15701 	(I27391,g27929);
	not 	XG15702 	(I26378,g26850);
	not 	XG15703 	(I26427,g26859);
	not 	XG15704 	(I26309,g26825);
	not 	XG15705 	(I27495,g27961);
	not 	XG15706 	(g29878,g28421);
	not 	XG15707 	(g29863,g28410);
	not 	XG15708 	(g29812,g28381);
	not 	XG15709 	(g29847,g28395);
	not 	XG15710 	(g29846,g28391);
	not 	XG15711 	(g29862,g28406);
	not 	XG15712 	(g29811,g28376);
	not 	XG15713 	(g29800,g28363);
	or 	XG15714 	(g32223,g29637,g31142);
	not 	XG15715 	(I26334,g26834);
	not 	XG15716 	(g29505,g29186);
	not 	XG15717 	(I26130,g26510);
	and 	XG15718 	(g30073,g28194,g1379);
	and 	XG15719 	(g29625,g14226,g28514);
	and 	XG15720 	(g29639,g11618,g28510);
	and 	XG15721 	(g27096,g16475,g26026);
	and 	XG15722 	(g27213,g16721,g26026);
	or 	XG15723 	(g28230,g14261,g27669);
	nand 	XG15724 	(I29314,I29313,g29501);
	not 	XG15725 	(g31658,I29242);
	not 	XG15726 	(g27187,I25882);
	not 	XG15727 	(g27163,I25869);
	or 	XG15728 	(g27126,g25787,g24378);
	and 	XG15729 	(g29567,g28593,g2357);
	and 	XG15730 	(g29974,g12914,g29173);
	and 	XG15731 	(g29988,g12235,g29187);
	and 	XG15732 	(g30071,g12975,g29184);
	and 	XG15733 	(g30082,g12752,g29181);
	and 	XG15734 	(g30070,g9529,g29167);
	and 	XG15735 	(g30060,g10581,g29146);
	and 	XG15736 	(g28283,g27445,g2361,g7380);
	or 	XG15737 	(g30279,g27668,g28637);
	and 	XG15738 	(g29350,g28395,g4939);
	not 	XG15739 	(g30012,I28241);
	and 	XG15740 	(g28799,g27445,g25348,g26424,g21434);
	and 	XG15741 	(g28761,g27416,g25299,g26424,g21434);
	and 	XG15742 	(g28833,g27469,g25388,g26424,g21434);
	and 	XG15743 	(g28789,g27440,g25340,g26424,g21434);
	and 	XG15744 	(g28739,g27395,g25274,g26424,g21434);
	and 	XG15745 	(g28846,g27474,g25399,g26424,g21434);
	and 	XG15746 	(g28768,g27421,g25308,g26424,g21434);
	and 	XG15747 	(g28880,g27494,g25438,g26424,g21434);
	nor 	XG15748 	(g29675,g8354,g8236,g28380);
	nor 	XG15749 	(g29705,g8404,g8284,g28399);
	and 	XG15750 	(g30007,g12929,g29141);
	and 	XG15751 	(g30027,g12550,g29104);
	and 	XG15752 	(g30006,g9259,g29032);
	and 	XG15753 	(g29989,g10489,g29006);
	and 	XG15754 	(g29575,g28604,g2066);
	not 	XG15755 	(g31616,I29214);
	nand 	XG15756 	(I29270,I29269,g29486);
	not 	XG15757 	(g31646,I29228);
	not 	XG15758 	(g31631,I29221);
	nand 	XG15759 	(I29285,I29284,g29489);
	or 	XG15760 	(g27405,g25968,g24572);
	and 	XG15761 	(g29565,g28590,g1932);
	or 	XG15762 	(g32247,g29686,g31168);
	and 	XG15763 	(g28267,g27421,g2227,g7328);
	and 	XG15764 	(g29578,g28606,g2491);
	and 	XG15765 	(g28291,g27469,g2070,g7411);
	and 	XG15766 	(g29632,g22417,g28899);
	and 	XG15767 	(g29523,g22417,g28930);
	and 	XG15768 	(g29533,g22417,g28958);
	and 	XG15769 	(g29991,g12922,g29179);
	and 	XG15770 	(g30008,g12297,g29191);
	and 	XG15771 	(g30033,g12937,g29189);
	and 	XG15772 	(g30045,g12419,g29200);
	and 	XG15773 	(g30032,g9326,g29072);
	and 	XG15774 	(g30015,g10519,g29040);
	and 	XG15775 	(g30029,g12936,g29164);
	and 	XG15776 	(g30042,g12601,g29142);
	or 	XG15777 	(g32211,g29603,g31124);
	and 	XG15778 	(g29536,g22432,g28969);
	and 	XG15779 	(g29614,g22369,g28860);
	and 	XG15780 	(g29516,g22369,g28895);
	and 	XG15781 	(g29569,g22498,g29028);
	and 	XG15782 	(g28293,g27474,g2495,g7424);
	not 	XG15783 	(g30301,I28548);
	or 	XG15784 	(g32218,g29619,g31130);
	not 	XG15785 	(g31624,I29218);
	not 	XG15786 	(g31639,I29225);
	nand 	XG15787 	(I29315,I29313,g12154);
	and 	XG15788 	(g29580,g14186,g28519);
	and 	XG15789 	(g29591,g11346,g28552);
	nand 	XG15790 	(I29286,I29284,g12085);
	not 	XG15791 	(I27449,g27737);
	and 	XG15792 	(g29611,g14209,g28540);
	and 	XG15793 	(g29626,g11415,g28584);
	and 	XG15794 	(g29610,g8026,g28483);
	and 	XG15795 	(g29595,g11833,g28475);
	or 	XG15796 	(g32264,g29711,g31187);
	and 	XG15797 	(g30011,g12930,g29183);
	and 	XG15798 	(g30030,g12347,g29198);
	and 	XG15799 	(g30010,g9274,g29035);
	and 	XG15800 	(g29992,g10490,g29012);
	and 	XG15801 	(g28439,g10233,g27273);
	and 	XG15802 	(g28254,g27395,g1668,g7268);
	and 	XG15803 	(g28889,g27395,g26424,g25169,g17292);
	not 	XG15804 	(g28918,g27832);
	and 	XG15805 	(g28924,g27416,g26424,g25183,g17317);
	and 	XG15806 	(g28281,g27440,g1936,g7362);
	and 	XG15807 	(g29607,g14208,g28509);
	and 	XG15808 	(g29623,g11563,g28496);
	nand 	XG15809 	(I29278,I29277,g29488);
	and 	XG15810 	(g29640,g8125,g28498);
	and 	XG15811 	(g29627,g11884,g28493);
	nand 	XG15812 	(I29279,I29277,g12081);
	nand 	XG15813 	(I29262,I29261,g29485);
	and 	XG15814 	(g30043,g9392,g29106);
	and 	XG15815 	(g30031,g10540,g29071);
	not 	XG15816 	(g29348,g28194);
	and 	XG15817 	(g29593,g7985,g28470);
	and 	XG15818 	(g29581,g11796,g28462);
	and 	XG15819 	(g30057,g9462,g29144);
	and 	XG15820 	(g30046,g10564,g29108);
	or 	XG15821 	(g30270,g27664,g28624);
	nand 	XG15822 	(g29355,g28109,g24383);
	nand 	XG15823 	(g29335,g28131,g25540);
	not 	XG15824 	(I28002,g28153);
	not 	XG15825 	(g30318,g28274);
	not 	XG15826 	(I28572,g28274);
	not 	XG15827 	(g29339,g28274);
	not 	XG15828 	(I28014,g28158);
	and 	XG15829 	(g31792,g24017,g30214);
	and 	XG15830 	(g31765,g23968,g30128);
	and 	XG15831 	(g31500,g23449,g29802);
	and 	XG15832 	(g31540,g23548,g29904);
	and 	XG15833 	(g29321,g22148,g29033);
	and 	XG15834 	(g31471,g23399,g29754);
	and 	XG15835 	(g31492,g23431,g29790);
	and 	XG15836 	(g31746,g23905,g30093);
	and 	XG15837 	(g31477,g23409,g29763);
	and 	XG15838 	(g29986,g23473,g28468);
	and 	XG15839 	(g31015,g22758,g29476);
	and 	XG15840 	(g31016,g22840,g29478);
	and 	XG15841 	(g31278,g23302,g29716);
	and 	XG15842 	(g31066,g22865,g29483);
	and 	XG15843 	(g31520,g23507,g29879);
	and 	XG15844 	(g31499,g23446,g29801);
	and 	XG15845 	(g31756,g23942,g30114);
	and 	XG15846 	(g31478,g23410,g29764);
	and 	XG15847 	(g29344,g18932,g29168);
	and 	XG15848 	(g31470,g23398,g29753);
	and 	XG15849 	(g31744,g23902,g30092);
	and 	XG15850 	(g32308,g23503,g31293);
	and 	XG15851 	(g31374,g23390,g29748);
	and 	XG15852 	(g30002,g23487,g28481);
	and 	XG15853 	(g31115,g22882,g29487);
	and 	XG15854 	(g31280,g23305,g29717);
	and 	XG15855 	(g31132,g22987,g29504);
	and 	XG15856 	(g31290,g23335,g29734);
	and 	XG15857 	(g31481,g23417,g29768);
	and 	XG15858 	(g32162,g23014,g31002);
	and 	XG15859 	(g31508,g23459,g29813);
	and 	XG15860 	(g31493,g23434,g29791);
	and 	XG15861 	(g31763,g23965,g30127);
	and 	XG15862 	(g31789,g24013,g30201);
	and 	XG15863 	(g31486,g23422,g29777);
	and 	XG15864 	(g31118,g22906,g29490);
	and 	XG15865 	(g31305,g23354,g29741);
	and 	XG15866 	(g31143,g22999,g29506);
	and 	XG15867 	(g31019,g22856,g29481);
	and 	XG15868 	(g27411,g17528,g26549);
	and 	XG15869 	(g27557,g17774,g26549);
	and 	XG15870 	(g27508,g17684,g26549);
	and 	XG15871 	(g27537,g17742,g26549);
	and 	XG15872 	(g27538,g14744,g26549);
	and 	XG15873 	(g27546,g17758,g26549);
	and 	XG15874 	(g27507,g17683,g26549);
	and 	XG15875 	(g27460,g17610,g26549);
	and 	XG15876 	(g27136,g16605,g26026);
	and 	XG15877 	(g27129,g16584,g26026);
	and 	XG15878 	(g27104,g16510,g25997);
	and 	XG15879 	(g27114,g16523,g25997);
	and 	XG15880 	(g27262,g17092,g25997);
	and 	XG15881 	(g27218,g16740,g25997);
	or 	XG15882 	(g27135,g25803,g24387);
	and 	XG15883 	(g27517,g17707,g26400);
	and 	XG15884 	(g27480,g17638,g26400);
	and 	XG15885 	(g27428,g17576,g26400);
	and 	XG15886 	(g27370,g17472,g26400);
	and 	XG15887 	(g27346,g17389,g26400);
	and 	XG15888 	(g27427,g17575,g26400);
	and 	XG15889 	(g27481,g14630,g26400);
	and 	XG15890 	(g27385,g17497,g26400);
	or 	XG15891 	(g32271,g29731,g31209);
	and 	XG15892 	(g27653,g15562,g26549);
	and 	XG15893 	(g27547,g17759,g26549);
	and 	XG15894 	(g27116,g16527,g26026);
	and 	XG15895 	(g27130,g16585,g26026);
	and 	XG15896 	(g27181,g16655,g26026);
	and 	XG15897 	(g27204,g16689,g26026);
	and 	XG15898 	(g29608,g11385,g28568);
	and 	XG15899 	(g29594,g14192,g28529);
	and 	XG15900 	(g30061,g28188,g1036);
	nand 	XG15901 	(I26438,g14271,g26549);
	and 	XG15902 	(g27220,g16743,g26026);
	and 	XG15903 	(g27203,g16688,g26026);
	and 	XG15904 	(g27106,g16512,g26026);
	and 	XG15905 	(g27151,g16626,g26026);
	and 	XG15906 	(g27115,g16526,g26026);
	and 	XG15907 	(g27214,g13901,g26026);
	and 	XG15908 	(g27219,g16742,g26026);
	and 	XG15909 	(g27137,g16606,g26026);
	and 	XG15910 	(g27105,g16511,g26026);
	and 	XG15911 	(g27180,g16654,g26026);
	and 	XG15912 	(g27373,g17477,g26488);
	and 	XG15913 	(g27387,g17499,g26488);
	and 	XG15914 	(g27267,g17124,g26026);
	and 	XG15915 	(g27227,g16771,g26026);
	not 	XG15916 	(I30904,g32424);
	and 	XG15917 	(g27134,g16602,g25997);
	and 	XG15918 	(g27177,g16651,g25997);
	and 	XG15919 	(g27103,g16509,g25997);
	and 	XG15920 	(g27095,g16473,g25997);
	and 	XG15921 	(g27212,g16717,g25997);
	and 	XG15922 	(g27211,g16716,g25997);
	and 	XG15923 	(g27094,g16472,g25997);
	and 	XG15924 	(g27202,g13876,g25997);
	and 	XG15925 	(g27148,g16622,g25997);
	and 	XG15926 	(g27128,g16583,g25997);
	and 	XG15927 	(g27645,g15344,g26488);
	and 	XG15928 	(g27534,g17735,g26488);
	and 	XG15929 	(g30050,g28126,g22545);
	not 	XG15930 	(g29342,g28188);
	and 	XG15931 	(g27389,g17503,g26519);
	and 	XG15932 	(g27486,g17645,g26519);
	and 	XG15933 	(g27545,g17756,g26519);
	and 	XG15934 	(g27520,g17714,g26519);
	and 	XG15935 	(g27521,g14700,g26519);
	and 	XG15936 	(g27433,g17583,g26519);
	and 	XG15937 	(g27485,g17644,g26519);
	and 	XG15938 	(g27535,g17737,g26519);
	and 	XG15939 	(g27650,g15479,g26519);
	and 	XG15940 	(g27536,g17738,g26519);
	and 	XG15941 	(g27347,g17390,g26400);
	and 	XG15942 	(g27371,g17473,g26400);
	and 	XG15943 	(g27500,g17672,g26400);
	and 	XG15944 	(g27358,g17415,g26400);
	and 	XG15945 	(g27437,g17589,g26576);
	and 	XG15946 	(g27462,g17612,g26576);
	or 	XG15947 	(g32243,g29683,g31166);
	nand 	XG15948 	(I29263,I29261,g12046);
	nand 	XG15949 	(I29296,I29295,g29495);
	and 	XG15950 	(g29552,g28579,g2223);
	or 	XG15951 	(g27431,g25977,g24582);
	and 	XG15952 	(g27207,g16692,g26055);
	and 	XG15953 	(g27132,g16589,g26055);
	and 	XG15954 	(g27234,g16814,g26055);
	and 	XG15955 	(g27221,g16747,g26055);
	and 	XG15956 	(g27206,g16691,g26055);
	and 	XG15957 	(g27154,g16630,g26055);
	and 	XG15958 	(g27228,g16773,g26055);
	and 	XG15959 	(g27222,g13932,g26055);
	and 	XG15960 	(g27272,g17144,g26055);
	and 	XG15961 	(g27229,g16774,g26055);
	nand 	XG15962 	(I29254,I29253,g29482);
	and 	XG15963 	(g27457,g17606,g26519);
	and 	XG15964 	(g27375,g17479,g26519);
	and 	XG15965 	(g27504,g17680,g26519);
	and 	XG15966 	(g27409,g17524,g26519);
	and 	XG15967 	(g27361,g17419,g26519);
	and 	XG15968 	(g27505,g17681,g26519);
	and 	XG15969 	(g27201,g16685,g25997);
	and 	XG15970 	(g27149,g16623,g25997);
	and 	XG15971 	(g27113,g16522,g25997);
	and 	XG15972 	(g27178,g16652,g25997);
	and 	XG15973 	(g27127,g16582,g25997);
	and 	XG15974 	(g27090,g16423,g25997);
	nand 	XG15975 	(I26070,g13517,g26026);
	and 	XG15976 	(g27372,g17476,g26488);
	and 	XG15977 	(g27360,g17417,g26488);
	and 	XG15978 	(g27482,g17641,g26488);
	and 	XG15979 	(g27430,g17579,g26488);
	and 	XG15980 	(g27519,g17710,g26488);
	and 	XG15981 	(g27518,g17709,g26488);
	and 	XG15982 	(g27454,g17602,g26488);
	and 	XG15983 	(g27407,g17522,g26488);
	and 	XG15984 	(g27359,g17416,g26488);
	and 	XG15985 	(g27503,g14668,g26488);
	and 	XG15986 	(g29590,g28615,g2625);
	and 	XG15987 	(g27490,g17651,g26576);
	and 	XG15988 	(g27461,g17611,g26576);
	and 	XG15989 	(g27526,g17721,g26576);
	and 	XG15990 	(g27540,g17746,g26576);
	and 	XG15991 	(g27215,g16724,g26055);
	and 	XG15992 	(g27183,g16658,g26055);
	and 	XG15993 	(g27118,g16529,g26055);
	and 	XG15994 	(g27216,g16725,g26055);
	and 	XG15995 	(g27139,g16608,g26055);
	and 	XG15996 	(g27107,g16514,g26055);
	and 	XG15997 	(g27404,g17518,g26400);
	and 	XG15998 	(g27357,g17414,g26400);
	and 	XG15999 	(g27501,g17673,g26400);
	and 	XG16000 	(g27451,g17599,g26400);
	and 	XG16001 	(g27628,g18061,g26400);
	and 	XG16002 	(g27339,g17308,g26400);
	and 	XG16003 	(g27452,g17600,g26400);
	and 	XG16004 	(g27384,g17496,g26400);
	nand 	XG16005 	(I26459,g14306,g26576);
	nand 	XG16006 	(I29255,I29253,g12017);
	or 	XG16007 	(g32210,g29600,g31123);
	and 	XG16008 	(g27376,g17481,g26549);
	and 	XG16009 	(g27522,g17717,g26549);
	and 	XG16010 	(g27390,g17504,g26549);
	and 	XG16011 	(g27410,g17527,g26549);
	and 	XG16012 	(g27434,g17584,g26549);
	and 	XG16013 	(g27459,g17609,g26549);
	or 	XG16014 	(g32285,g29740,g31222);
	or 	XG16015 	(g32229,g29652,g31148);
	and 	XG16016 	(g27408,g17523,g26519);
	and 	XG16017 	(g27374,g17478,g26519);
	and 	XG16018 	(g27432,g17582,g26519);
	and 	XG16019 	(g27388,g17502,g26519);
	nand 	XG16020 	(I29271,I29269,g12050);
	and 	XG16021 	(g27117,g16528,g26055);
	and 	XG16022 	(g27131,g16588,g26055);
	and 	XG16023 	(g27138,g16607,g26055);
	and 	XG16024 	(g27153,g16629,g26055);
	not 	XG16025 	(g28754,I27238);
	or 	XG16026 	(g32216,g29615,g31128);
	nand 	XG16027 	(I26366,g14211,g26400);
	nand 	XG16028 	(I26049,g13500,g25997);
	and 	XG16029 	(g27455,g17603,g26488);
	and 	XG16030 	(g27386,g17498,g26488);
	and 	XG16031 	(g27502,g17677,g26488);
	and 	XG16032 	(g27348,g17392,g26488);
	and 	XG16033 	(g27483,g17642,g26488);
	and 	XG16034 	(g27406,g17521,g26488);
	and 	XG16035 	(g27391,g17505,g26549);
	and 	XG16036 	(g27488,g17648,g26549);
	and 	XG16037 	(g27435,g17585,g26549);
	and 	XG16038 	(g27523,g17718,g26549);
	nand 	XG16039 	(I26393,g14227,g26488);
	or 	XG16040 	(g32277,g29733,g31211);
	and 	XG16041 	(g29537,g22472,g28976);
	and 	XG16042 	(g29618,g22384,g28870);
	and 	XG16043 	(g29518,g22384,g28906);
	nand 	XG16044 	(I29303,I29302,g29496);
	and 	XG16045 	(g27525,g17720,g26576);
	and 	XG16046 	(g27412,g17529,g26576);
	and 	XG16047 	(g27558,g17776,g26576);
	and 	XG16048 	(g27549,g14785,g26576);
	and 	XG16049 	(g27491,g17652,g26576);
	and 	XG16050 	(g27436,g17588,g26576);
	and 	XG16051 	(g27413,g17530,g26576);
	and 	XG16052 	(g27539,g17745,g26576);
	and 	XG16053 	(g27559,g17777,g26576);
	and 	XG16054 	(g27510,g17687,g26576);
	or 	XG16055 	(g32237,g29667,g31153);
	or 	XG16056 	(g32235,g29662,g31151);
	nand 	XG16057 	(I29304,I29302,g12121);
	nand 	XG16058 	(I26417,g14247,g26519);
	and 	XG16059 	(g27548,g17763,g26576);
	and 	XG16060 	(g27568,g17791,g26576);
	and 	XG16061 	(g27392,g17507,g26576);
	and 	XG16062 	(g27661,g15568,g26576);
	nand 	XG16063 	(I26093,g13539,g26055);
	or 	XG16064 	(g32259,g29709,g31185);
	nand 	XG16065 	(I29297,I29295,g12117);
	or 	XG16066 	(g27383,g25961,g24569);
	or 	XG16067 	(g32976,g21704,g32207);
	or 	XG16068 	(g32209,g29599,g31122);
	or 	XG16069 	(g32233,g29661,g31150);
	or 	XG16070 	(g32220,g29633,g31139);
	or 	XG16071 	(g32221,g29634,g31140);
	and 	XG16072 	(g29526,g22384,g28938);
	and 	XG16073 	(g29650,g22472,g28949);
	and 	XG16074 	(g29554,g22472,g28997);
	or 	XG16075 	(g32217,g29616,g31129);
	and 	XG16076 	(g29527,g22432,g28945);
	and 	XG16077 	(g29635,g22432,g28910);
	and 	XG16078 	(g29666,g22498,g28980);
	and 	XG16079 	(g29555,g22498,g29004);
	or 	XG16080 	(g32227,g29648,g31146);
	or 	XG16081 	(g32982,g18208,g31948);
	or 	XG16082 	(g32981,g18206,g32425);
	and 	XG16083 	(g33723,g33299,g14091);
	nor 	XG16084 	(g33851,g12259,g33299,g8854);
	or 	XG16085 	(g32977,g21710,g32169);
	or 	XG16086 	(g27152,g25817,g24393);
	or 	XG16087 	(g32208,g29584,g31120);
	not 	XG16088 	(g31795,I29371);
	not 	XG16089 	(I29717,g30931);
	not 	XG16090 	(I29720,g30931);
	and 	XG16091 	(g30035,g28120,g22539);
	or 	XG16092 	(g33123,g30577,g31962);
	or 	XG16093 	(g32980,g18198,g32254);
	not 	XG16094 	(g33799,g33299);
	or 	XG16095 	(g32226,g29645,g31145);
	and 	XG16096 	(g33102,g18978,g32399);
	and 	XG16097 	(g33099,g18944,g32395);
	and 	XG16098 	(g33817,g20102,g33235);
	and 	XG16099 	(g33186,g22830,g32037);
	and 	XG16100 	(g33241,g23128,g32173);
	and 	XG16101 	(g33245,g19961,g32125);
	and 	XG16102 	(g33122,g32192,g8859);
	or 	XG16103 	(g33232,g30936,g32034);
	and 	XG16104 	(g33724,g33258,g14145);
	or 	XG16105 	(g27458,g25989,g24590);
	or 	XG16106 	(g33615,g21871,g33113);
	or 	XG16107 	(g32257,g29708,g31184);
	or 	XG16108 	(g27489,g26022,g24608);
	or 	XG16109 	(g33794,g32053,g33126);
	or 	XG16110 	(g32245,g29684,g31167);
	or 	XG16111 	(g27159,g12953,g25814);
	or 	XG16112 	(g32985,g18266,g31963);
	or 	XG16113 	(g31872,g18535,g31524);
	or 	XG16114 	(g33019,g18536,g32339);
	and 	XG16115 	(g33121,g32212,g8748);
	nand 	XG16116 	(g33306,g11679,g32212,g776);
	and 	XG16117 	(g33104,g32137,g26296);
	or 	XG16118 	(g32984,g18264,g31934);
	or 	XG16119 	(g33291,g13477,g32154);
	and 	XG16120 	(g33244,g23152,g32190);
	or 	XG16121 	(g33538,g18144,g33252);
	and 	XG16122 	(g33233,g23005,g32094);
	not 	XG16123 	(g33246,g32212);
	or 	XG16124 	(g32979,g18177,g32181);
	and 	XG16125 	(g33322,g20450,g32202);
	and 	XG16126 	(g33105,g32138,g26298);
	or 	XG16127 	(g33159,g30730,g32016);
	not 	XG16128 	(g30326,I28579);
	not 	XG16129 	(g28436,I26929);
	not 	XG16130 	(g28463,I26952);
	and 	XG16131 	(g29752,g10233,g28516);
	and 	XG16132 	(g29736,g10233,g28522);
	and 	XG16133 	(g29718,g11136,g28512);
	not 	XG16134 	(I28480,g28652);
	not 	XG16135 	(g27438,I26130);
	and 	XG16136 	(g30599,g29863,g18911);
	and 	XG16137 	(g30595,g29847,g18911);
	and 	XG16138 	(g30604,g29878,g18911);
	and 	XG16139 	(g30590,g29812,g18911);
	not 	XG16140 	(I29204,g29505);
	or 	XG16141 	(g31248,g29522,g25970);
	or 	XG16142 	(g31241,g29510,g25959);
	or 	XG16143 	(g31257,g28253,g29531);
	not 	XG16144 	(g27708,I26334);
	or 	XG16145 	(g31258,g29550,g25991);
	or 	XG16146 	(g31254,g29534,g25981);
	and 	XG16147 	(g29966,g28970,g23617);
	and 	XG16148 	(g31376,g29814,g24952);
	and 	XG16149 	(g30735,g22319,g29814);
	and 	XG16150 	(g31514,g29956,g20041);
	and 	XG16151 	(g31497,g29930,g20041);
	and 	XG16152 	(g31503,g29945,g20041);
	and 	XG16153 	(g31518,g29970,g20041);
	or 	XG16154 	(g33066,g22096,g32341);
	and 	XG16155 	(g32126,g29948,g31601);
	and 	XG16156 	(g32106,g29911,g31601);
	not 	XG16157 	(g29195,I27495);
	and 	XG16158 	(g31223,g29689,g20028);
	and 	XG16159 	(g31212,g29669,g20028);
	and 	XG16160 	(g31228,g29713,g20028);
	and 	XG16161 	(g31188,g29653,g20028);
	or 	XG16162 	(g30457,g21885,g29369);
	not 	XG16163 	(g27675,I26309);
	or 	XG16164 	(g30459,g21926,g29314);
	or 	XG16165 	(g31465,g29647,g26156);
	or 	XG16166 	(g31295,g29598,g26090);
	not 	XG16167 	(g27880,I26427);
	and 	XG16168 	(g32234,g30292,g31601);
	and 	XG16169 	(g32096,g29893,g31601);
	or 	XG16170 	(g31919,g22044,g31758);
	and 	XG16171 	(g29952,g28939,g23576);
	not 	XG16172 	(g27773,I26378);
	or 	XG16173 	(g31267,g28263,g29548);
	not 	XG16174 	(g29043,I27391);
	not 	XG16175 	(g27709,I26337);
	and 	XG16176 	(g29979,g28991,g23655);
	not 	XG16177 	(I26880,g27527);
	or 	XG16178 	(I28567,g29207,g29206,g29205,g29204);
	or 	XG16179 	(I28566,g28035,g29203,g29202,g29201);
	or 	XG16180 	(g28220,I26742,I26741,g23495);
	or 	XG16181 	(g31931,g22095,g31494);
	not 	XG16182 	(g27013,I25743);
	not 	XG16183 	(g30997,g29702);
	not 	XG16184 	(g30999,g29722);
	and 	XG16185 	(g29982,g28998,g23656);
	or 	XG16186 	(g29529,g28267,g28283,g28293,g28303);
	not 	XG16187 	(g29013,I27368);
	not 	XG16188 	(I27314,g28009);
	or 	XG16189 	(g31928,g22092,g31517);
	not 	XG16190 	(g30989,g29672);
	not 	XG16191 	(g30996,g29694);
	not 	XG16192 	(g30990,g29676);
	not 	XG16193 	(g31000,g29737);
	not 	XG16194 	(I28851,g29317);
	not 	XG16195 	(g27998,I26512);
	nand 	XG16196 	(g31003,g19644,g29497,g27163);
	nand 	XG16197 	(g31009,g19644,g29503,g27187);
	or 	XG16198 	(g30337,g18220,g29334);
	not 	XG16199 	(g30217,I28458);
	or 	XG16200 	(g31888,g21821,g31067);
	and 	XG16201 	(g29810,g11317,g28259);
	and 	XG16202 	(g29789,g10233,g28270);
	and 	XG16203 	(g29773,g10233,g28203);
	and 	XG16204 	(g29762,g10233,g28298);
	and 	XG16205 	(g29743,g10233,g28206);
	and 	XG16206 	(g29742,g10233,g28288);
	and 	XG16207 	(g29774,g10233,g28287);
	and 	XG16208 	(g29693,g10233,g28207);
	and 	XG16209 	(g29799,g10233,g28271);
	or 	XG16210 	(g31922,g22047,g31525);
	or 	XG16211 	(g31901,g21909,g31516);
	or 	XG16212 	(g31913,g21999,g31485);
	not 	XG16213 	(g27736,I26356);
	and 	XG16214 	(g32139,g29960,g31601);
	and 	XG16215 	(g32113,g29925,g31601);
	or 	XG16216 	(g33051,g21958,g32316);
	and 	XG16217 	(g29962,g28959,g23616);
	or 	XG16218 	(g29520,g28254,g28264,g28281,g28291);
	or 	XG16219 	(g31885,g21779,g31017);
	or 	XG16220 	(g31775,g30059,g30048);
	not 	XG16221 	(I27253,g27996);
	or 	XG16222 	(g31911,g21969,g31784);
	and 	XG16223 	(g31070,g25985,g29814);
	and 	XG16224 	(g30937,g29814,g22626);
	and 	XG16225 	(g31021,g29814,g26025);
	and 	XG16226 	(g31554,g29814,g19050);
	and 	XG16227 	(g31566,g29814,g19050);
	and 	XG16228 	(g31528,g29814,g19050);
	and 	XG16229 	(g31672,g19050,g29814);
	and 	XG16230 	(g31542,g29814,g19050);
	and 	XG16231 	(g31579,g29814,g19128);
	and 	XG16232 	(g31710,g19128,g29814);
	and 	XG16233 	(g31170,g29814,g19128);
	and 	XG16234 	(g31194,g29814,g19128);
	and 	XG16235 	(g31154,g29814,g19128);
	and 	XG16236 	(g31327,g29814,g19200);
	or 	XG16237 	(g30435,g21840,g30025);
	or 	XG16238 	(g31876,g21731,g31125);
	or 	XG16239 	(g31908,g21955,g31519);
	and 	XG16240 	(g30000,g29029,g23685);
	and 	XG16241 	(g32140,g29961,g31609);
	and 	XG16242 	(g32109,g29920,g31609);
	not 	XG16243 	(I27232,g27993);
	not 	XG16244 	(g27967,I26479);
	or 	XG16245 	(g31893,g21837,g31490);
	or 	XG16246 	(g31468,g29656,g29641);
	not 	XG16247 	(I27738,g28140);
	or 	XG16248 	(g30501,g22018,g29327);
	not 	XG16249 	(I27388,g27698);
	or 	XG16250 	(g31904,g21923,g31780);
	not 	XG16251 	(g30983,g29657);
	not 	XG16252 	(g30998,g29719);
	or 	XG16253 	(g31770,g30047,g30034);
	or 	XG16254 	(g31745,g29973,g29959);
	or 	XG16255 	(g31887,g21820,g31292);
	or 	XG16256 	(g31918,g22015,g31786);
	or 	XG16257 	(g31773,g30056,g30044);
	or 	XG16258 	(g31900,g21908,g31484);
	or 	XG16259 	(g33030,g21826,g32166);
	not 	XG16260 	(g29311,g28998);
	not 	XG16261 	(g29318,g29029);
	or 	XG16262 	(g31898,g21906,g31707);
	not 	XG16263 	(g27774,I26381);
	and 	XG16264 	(g30614,g29814,g20154);
	and 	XG16265 	(g30825,g22332,g29814);
	and 	XG16266 	(g30673,g29814,g20175);
	or 	XG16267 	(g31912,g21998,g31752);
	or 	XG16268 	(g33056,g22004,g32327);
	not 	XG16269 	(I29337,g30286);
	not 	XG16270 	(g30309,g28959);
	not 	XG16271 	(g29310,g28991);
	or 	XG16272 	(g31761,g30028,g30009);
	or 	XG16273 	(g30543,g22110,g29338);
	or 	XG16274 	(g31316,g29624,g29609);
	or 	XG16275 	(g31751,g29990,g29975);
	or 	XG16276 	(g31930,g22094,g31769);
	or 	XG16277 	(g31881,g21775,g31018);
	or 	XG16278 	(g31873,g21728,g31270);
	or 	XG16279 	(g31909,g21956,g31750);
	or 	XG16280 	(g33020,g21734,g32160);
	not 	XG16281 	(g30305,g28939);
	not 	XG16282 	(g30312,g28970);
	not 	XG16283 	(g27928,g26810);
	or 	XG16284 	(g30522,g22064,g29332);
	not 	XG16285 	(g27930,I26451);
	not 	XG16286 	(g27956,I26466);
	or 	XG16287 	(g31781,g30069,g30058);
	or 	XG16288 	(g33061,g22050,g32334);
	not 	XG16289 	(g27830,g26802);
	or 	XG16290 	(g31303,g29606,g29592);
	or 	XG16291 	(g31279,g29579,g29571);
	or 	XG16292 	(g31879,g21745,g31475);
	nor 	XG16293 	(g30934,g29850,g29836);
	nor 	XG16294 	(g30929,g29835,g29803);
	nor 	XG16295 	(g31008,g30026,g30004);
	not 	XG16296 	(g30195,I28434);
	not 	XG16297 	(g29365,g29067);
	not 	XG16298 	(g30578,g29956);
	not 	XG16299 	(g30593,g29970);
	not 	XG16300 	(g31608,g29653);
	not 	XG16301 	(g30572,g29945);
	not 	XG16302 	(g31623,g29669);
	not 	XG16303 	(g31638,g29689);
	not 	XG16304 	(g31653,g29713);
	not 	XG16305 	(g30567,g29930);
	and 	XG16306 	(g33344,g20670,g32228);
	and 	XG16307 	(g33341,g20640,g32223);
	and 	XG16308 	(g33364,g20921,g32264);
	and 	XG16309 	(g33368,g21057,g32275);
	and 	XG16310 	(g28542,g20275,g27405);
	and 	XG16311 	(g33340,g20639,g32222);
	and 	XG16312 	(g33358,g20778,g32249);
	and 	XG16313 	(g33363,g20918,g32262);
	and 	XG16314 	(g33334,g20613,g32219);
	and 	XG16315 	(g28228,g19636,g27126);
	and 	XG16316 	(g33357,g20775,g32247);
	and 	XG16317 	(g33330,g20588,g32211);
	and 	XG16318 	(g33333,g20612,g32218);
	and 	XG16319 	(g33351,g20707,g32236);
	and 	XG16320 	(g30005,g24394,g28230);
	and 	XG16321 	(g30596,g18947,g30279);
	and 	XG16322 	(g30592,g18929,g30270);
	and 	XG16323 	(g28224,g27064,g22763,g27163);
	not 	XG16324 	(g29765,I28014);
	not 	XG16325 	(g30568,g29339);
	not 	XG16326 	(g30321,I28572);
	and 	XG16327 	(g29382,g28172,g22763,g26424);
	not 	XG16328 	(g29755,I28002);
	and 	XG16329 	(g28231,g27074,g22763,g27187);
	and 	XG16330 	(g29384,g28179,g22763,g26424);
	and 	XG16331 	(g32119,g29939,g31609);
	and 	XG16332 	(g32145,g29977,g31609);
	and 	XG16333 	(g29949,g28924,g23575);
	or 	XG16334 	(g29366,g28439,g13738);
	or 	XG16335 	(g29373,g28453,g13832);
	or 	XG16336 	(g31253,g29533,g25980);
	or 	XG16337 	(g31774,g30057,g30046);
	and 	XG16338 	(g32127,g29950,g31624);
	and 	XG16339 	(g32107,g29912,g31624);
	nor 	XG16340 	(g30156,g14587,g28789);
	nor 	XG16341 	(g30144,g7322,g28789);
	nor 	XG16342 	(g32017,g23475,g31504);
	or 	XG16343 	(g31291,g29593,g29581);
	or 	XG16344 	(g31274,g28280,g29565);
	or 	XG16345 	(g31249,g29523,g25971);
	and 	XG16346 	(g32108,g29913,g31631);
	nor 	XG16347 	(g30159,g14589,g28799);
	and 	XG16348 	(g32128,g29953,g31631);
	nor 	XG16349 	(g30148,g7335,g28799);
	and 	XG16350 	(g32122,g29944,g31646);
	and 	XG16351 	(g32153,g29999,g31646);
	nor 	XG16352 	(g30150,g7424,g28846);
	and 	XG16353 	(g32103,g29905,g31609);
	nor 	XG16354 	(g30143,g14566,g28761);
	and 	XG16355 	(g32244,g30297,g31609);
	nor 	XG16356 	(g30130,g7275,g28761);
	or 	XG16357 	(g31276,g28282,g29567);
	or 	XG16358 	(g28297,g15785,g27096);
	or 	XG16359 	(g31767,g30043,g30031);
	and 	XG16360 	(g32129,g29955,g31658);
	and 	XG16361 	(g32158,g30022,g31658);
	nor 	XG16362 	(g30162,g7462,g28880);
	and 	XG16363 	(g28141,g27163,g11261,g11797,g10831);
	and 	XG16364 	(g30576,g29800,g18898);
	and 	XG16365 	(g30594,g29846,g18898);
	and 	XG16366 	(g30589,g29811,g18898);
	and 	XG16367 	(g30598,g29862,g18898);
	nand 	XG16368 	(g31671,I29263,I29262);
	nand 	XG16369 	(g31708,I29279,I29278);
	or 	XG16370 	(g31326,g29640,g29627);
	nor 	XG16371 	(g30119,g7315,g28761);
	and 	XG16372 	(g32149,g29983,g31658);
	and 	XG16373 	(g32159,g30040,g31658);
	nor 	XG16374 	(g30183,g14644,g28880);
	or 	XG16375 	(g31315,g29623,g29607);
	or 	XG16376 	(g31308,g29614,g26101);
	or 	XG16377 	(g31269,g29569,g26024);
	and 	XG16378 	(g32150,g29995,g31624);
	and 	XG16379 	(g32258,g30303,g31624);
	not 	XG16380 	(g30302,g28924);
	not 	XG16381 	(g30218,g28918);
	not 	XG16382 	(g30296,g28889);
	and 	XG16383 	(g32151,g29996,g31639);
	and 	XG16384 	(g32120,g29941,g31639);
	nor 	XG16385 	(g30146,g7411,g28833);
	or 	XG16386 	(g31255,g29536,g25982);
	or 	XG16387 	(g31320,g29632,g26125);
	and 	XG16388 	(g32116,g29929,g31658);
	and 	XG16389 	(g32286,g29312,g31658);
	nor 	XG16390 	(g30171,g7431,g28880);
	or 	XG16391 	(g31757,g30010,g29992);
	or 	XG16392 	(g31762,g30030,g30011);
	and 	XG16393 	(g32114,g29927,g31624);
	and 	XG16394 	(g32146,g29978,g31624);
	nor 	XG16395 	(g30132,g7362,g28789);
	nand 	XG16396 	(g31706,I29271,I29270);
	and 	XG16397 	(g32104,g29906,g31616);
	nor 	XG16398 	(g30147,g14567,g28768);
	and 	XG16399 	(g32121,g29942,g31616);
	nor 	XG16400 	(g30134,g7280,g28768);
	or 	XG16401 	(g31306,g29610,g29595);
	or 	XG16402 	(g31317,g29626,g29611);
	or 	XG16403 	(g31287,g28292,g29578);
	not 	XG16404 	(g29147,I27449);
	or 	XG16405 	(g31244,g29515,g25963);
	nand 	XG16406 	(g31709,I29286,I29285);
	nand 	XG16407 	(g28336,g19644,g27163,g24756,g27064);
	nand 	XG16408 	(g28349,g19644,g27187,g24770,g27074);
	or 	XG16409 	(g31289,g29591,g29580);
	nand 	XG16410 	(g31753,I29315,I29314);
	not 	XG16411 	(I28832,g30301);
	and 	XG16412 	(g28150,g27187,g11283,g11834,g10862);
	and 	XG16413 	(g32157,g30021,g31646);
	and 	XG16414 	(g32143,g29967,g31646);
	nor 	XG16415 	(g30170,g14615,g28846);
	or 	XG16416 	(g31766,g30042,g30029);
	or 	XG16417 	(g31764,g30032,g30015);
	or 	XG16418 	(g31768,g30045,g30033);
	or 	XG16419 	(g31755,g30008,g29991);
	nor 	XG16420 	(g30169,g14613,g28833);
	and 	XG16421 	(g32148,g29981,g31631);
	and 	XG16422 	(g32115,g29928,g31631);
	nor 	XG16423 	(g30136,g7380,g28799);
	and 	XG16424 	(g32147,g29980,g31616);
	and 	XG16425 	(g32248,g30299,g31616);
	nor 	XG16426 	(g30129,g14537,g28739);
	nor 	XG16427 	(g30117,g7252,g28739);
	or 	XG16428 	(g31284,g28290,g29575);
	or 	XG16429 	(g31754,g30006,g29989);
	or 	XG16430 	(g31760,g30027,g30007);
	not 	XG16431 	(I29013,g29705);
	not 	XG16432 	(I29002,g29675);
	nor 	XG16433 	(g30106,g7268,g28739);
	nor 	XG16434 	(g30123,g7328,g28768);
	nor 	XG16435 	(g30160,g7387,g28846);
	and 	XG16436 	(g28484,I26972,g21163,g10290,g27187);
	and 	XG16437 	(g29073,I27409,g21012,g10290,g27163);
	and 	XG16438 	(g29192,g10290,g27163);
	and 	XG16439 	(g28553,g10290,g27187);
	and 	XG16440 	(g29182,g12730,g27163);
	and 	XG16441 	(g29008,I27364,g20739,g12730,g27163);
	and 	XG16442 	(g28528,g12730,g27187);
	and 	XG16443 	(g28458,I26948,g20887,g12730,g27187);
	not 	XG16444 	(I29185,g30012);
	not 	XG16445 	(I29182,g30012);
	or 	XG16446 	(g28402,g15873,g27213);
	or 	XG16447 	(g31782,g30070,g30060);
	or 	XG16448 	(g31785,g30082,g30071);
	or 	XG16449 	(g31749,g29988,g29974);
	and 	XG16450 	(g28471,I26960,g21024,g12762,g27187);
	and 	XG16451 	(g29036,I27381,g20875,g12762,g27163);
	and 	XG16452 	(g29188,g12762,g27163);
	and 	XG16453 	(g28539,g12762,g27187);
	and 	XG16454 	(g29199,g12687,g27187);
	and 	XG16455 	(g28982,I27349,g20682,g12687,g27163);
	and 	XG16456 	(g29178,g12687,g27163);
	and 	XG16457 	(g29110,I27429,g20751,g12687,g27187);
	or 	XG16458 	(g29197,g27163,g27187);
	or 	XG16459 	(g31325,g29639,g29625);
	or 	XG16460 	(g29105,g17134,g27645);
	and 	XG16461 	(g31541,g29348,g22536);
	nor 	XG16462 	(g30157,g7369,g28833);
	and 	XG16463 	(g32272,g30310,g31639);
	and 	XG16464 	(g32110,g29921,g31639);
	or 	XG16465 	(g28342,g15819,g27134);
	or 	XG16466 	(g28659,g16610,g27404);
	or 	XG16467 	(g28316,g15804,g27113);
	or 	XG16468 	(g31905,g21952,g31746);
	or 	XG16469 	(g33025,g21780,g32162);
	or 	XG16470 	(g28371,g15847,g27177);
	nand 	XG16471 	(I26094,I26093,g26055);
	nand 	XG16472 	(I26367,I26366,g26400);
	nand 	XG16473 	(I26050,I26049,g25997);
	nand 	XG16474 	(I26394,I26393,g26488);
	nand 	XG16475 	(I26418,I26417,g26519);
	nand 	XG16476 	(I26460,I26459,g26576);
	nand 	XG16477 	(I26071,I26070,g26026);
	nand 	XG16478 	(I26439,I26438,g26549);
	or 	XG16479 	(g28357,g15836,g27148);
	nand 	XG16480 	(g31747,I29297,I29296);
	or 	XG16481 	(g28705,g16672,g27460);
	or 	XG16482 	(g29068,g17119,g27628);
	or 	XG16483 	(g28497,g16199,g27267);
	or 	XG16484 	(g28632,g16535,g27373);
	or 	XG16485 	(g28416,g15880,g27218);
	or 	XG16486 	(g28404,g15874,g27215);
	or 	XG16487 	(g29176,g17177,g27661);
	or 	XG16488 	(g31902,g21910,g31744);
	or 	XG16489 	(g31903,g21911,g31374);
	or 	XG16490 	(g28698,g16666,g27451);
	or 	XG16491 	(g31924,g22049,g31486);
	or 	XG16492 	(g28375,g15851,g27183);
	or 	XG16493 	(g31889,g21822,g31118);
	or 	XG16494 	(g28721,g16705,g27488);
	or 	XG16495 	(g28644,g16593,g27387);
	or 	XG16496 	(g28707,g16673,g27461);
	or 	XG16497 	(g28731,g16733,g27504);
	or 	XG16498 	(g28358,g15837,g27149);
	or 	XG16499 	(g31926,g22090,g31765);
	or 	XG16500 	(g28435,g15967,g27234);
	or 	XG16501 	(g28386,g13277,g27202);
	or 	XG16502 	(g28702,g16670,g27457);
	or 	XG16503 	(g31914,g22000,g31499);
	or 	XG16504 	(g28332,g15815,g27130);
	and 	XG16505 	(g32263,g30306,g31631);
	and 	XG16506 	(g32152,g29998,g31631);
	or 	XG16507 	(g28295,g15783,g27094);
	or 	XG16508 	(g28619,g16517,g27358);
	or 	XG16509 	(g28372,g15848,g27178);
	or 	XG16510 	(g28286,g15757,g27090);
	or 	XG16511 	(g28814,g16841,g27545);
	or 	XG16512 	(g28385,g15857,g27201);
	or 	XG16513 	(g31899,g21907,g31470);
	or 	XG16514 	(g28618,g16516,g27357);
	or 	XG16515 	(g28388,g15859,g27204);
	or 	XG16516 	(g28852,g16871,g27559);
	or 	XG16517 	(g28750,g16765,g27525);
	or 	XG16518 	(g31882,g21776,g31115);
	or 	XG16519 	(g28651,g16599,g27392);
	or 	XG16520 	(g28305,g15793,g27103);
	or 	XG16521 	(g28335,g15818,g27132);
	or 	XG16522 	(g30343,g18278,g29344);
	and 	XG16523 	(g32276,g30313,g31646);
	and 	XG16524 	(g32112,g29923,g31646);
	and 	XG16525 	(g32111,g29922,g31616);
	and 	XG16526 	(g32142,g29965,g31616);
	nand 	XG16527 	(I26419,I26417,g14247);
	or 	XG16528 	(g31906,g21953,g31477);
	or 	XG16529 	(g28334,g15817,g27131);
	or 	XG16530 	(g28734,g16736,g27508);
	or 	XG16531 	(g28691,g16642,g27437);
	nand 	XG16532 	(g31748,I29304,I29303);
	or 	XG16533 	(g31929,g22093,g31540);
	or 	XG16534 	(g28629,g16532,g27371);
	or 	XG16535 	(g28647,g16596,g27389);
	or 	XG16536 	(g31890,g21823,g31143);
	or 	XG16537 	(g30393,g21748,g29986);
	or 	XG16538 	(g28646,g16595,g27388);
	or 	XG16539 	(g31932,g22107,g31792);
	or 	XG16540 	(g28320,g15808,g27116);
	or 	XG16541 	(g28728,g16730,g27501);
	or 	XG16542 	(g31245,g29516,g25964);
	or 	XG16543 	(g31915,g22001,g31520);
	or 	XG16544 	(g28348,g15823,g27139);
	or 	XG16545 	(g28649,g16597,g27390);
	or 	XG16546 	(g28611,g16485,g27348);
	and 	XG16547 	(g32141,g29963,g31639);
	and 	XG16548 	(g32156,g30018,g31639);
	or 	XG16549 	(g31311,g29618,g26103);
	or 	XG16550 	(g28347,g15822,g27138);
	or 	XG16551 	(g28640,g16590,g27384);
	or 	XG16552 	(g28403,g13282,g27214);
	or 	XG16553 	(g31877,g21732,g31278);
	and 	XG16554 	(g30583,g29355,g19666);
	nand 	XG16555 	(g30573,g19666,g29355);
	nand 	XG16556 	(g30580,g19666,g29335);
	or 	XG16557 	(g28610,g16484,g27347);
	or 	XG16558 	(g28665,g16614,g27409);
	or 	XG16559 	(g28362,g15840,g27154);
	or 	XG16560 	(g28775,g16806,g27537);
	or 	XG16561 	(g28717,g16701,g27482);
	or 	XG16562 	(g28609,g16483,g27346);
	or 	XG16563 	(g28664,g16613,g27408);
	nand 	XG16564 	(I26395,I26393,g14227);
	or 	XG16565 	(g28361,g15839,g27153);
	or 	XG16566 	(g31927,g22091,g31500);
	or 	XG16567 	(g31268,g28266,g29552);
	or 	XG16568 	(g28662,g16612,g27407);
	or 	XG16569 	(g28685,g16637,g27433);
	or 	XG16570 	(g28323,g15810,g27118);
	or 	XG16571 	(g28684,g16636,g27432);
	or 	XG16572 	(g31923,g22048,g31763);
	or 	XG16573 	(g31878,g21733,g31015);
	or 	XG16574 	(g31910,g21957,g31471);
	or 	XG16575 	(g28635,g16537,g27375);
	or 	XG16576 	(g31880,g21774,g31280);
	not 	XG16577 	(g30142,g28754);
	or 	XG16578 	(g28778,g16808,g27540);
	or 	XG16579 	(g28727,g16729,g27500);
	or 	XG16580 	(g31886,g21791,g31481);
	or 	XG16581 	(g28743,g16758,g27517);
	or 	XG16582 	(g28428,g15912,g27227);
	or 	XG16583 	(g28490,g16185,g27262);
	or 	XG16584 	(g31874,g21729,g31016);
	or 	XG16585 	(g28373,g15849,g27180);
	or 	XG16586 	(g28329,g15813,g27128);
	or 	XG16587 	(g31907,g21954,g31492);
	or 	XG16588 	(g28641,g16591,g27385);
	and 	XG16589 	(g29938,g28889,g23552);
	nand 	XG16590 	(g31669,I29255,I29254);
	or 	XG16591 	(g28401,g15871,g27212);
	nand 	XG16592 	(I26461,I26459,g14306);
	or 	XG16593 	(g28328,g15812,g27127);
	or 	XG16594 	(g28680,g16633,g27427);
	or 	XG16595 	(g28417,g15881,g27219);
	or 	XG16596 	(g28344,g15820,g27136);
	or 	XG16597 	(g28621,g16518,g27359);
	or 	XG16598 	(g28359,g15838,g27151);
	or 	XG16599 	(g28600,g16427,g27339);
	or 	XG16600 	(g31875,g21730,g31066);
	or 	XG16601 	(g28420,g13290,g27222);
	or 	XG16602 	(g28723,g16706,g27490);
	or 	XG16603 	(g31302,g28302,g29590);
	or 	XG16604 	(g28733,g16735,g27507);
	or 	XG16605 	(g30480,g21972,g29321);
	or 	XG16606 	(g28390,g15861,g27207);
	or 	XG16607 	(g28747,g13942,g27521);
	or 	XG16608 	(g31891,g21824,g31305);
	or 	XG16609 	(g33046,g21912,g32308);
	or 	XG16610 	(g29166,g17153,g27653);
	or 	XG16611 	(g28720,g16704,g27486);
	or 	XG16612 	(g31916,g22002,g31756);
	or 	XG16613 	(g28815,g16842,g27546);
	or 	XG16614 	(g28715,g16700,g27480);
	or 	XG16615 	(g28400,g15870,g27211);
	or 	XG16616 	(g28776,g13974,g27538);
	or 	XG16617 	(g31892,g21825,g31019);
	or 	XG16618 	(g28331,g15814,g27129);
	or 	XG16619 	(g31779,g28673,g30050);
	or 	XG16620 	(g28816,g16843,g27547);
	not 	XG16621 	(g33378,I30904);
	or 	XG16622 	(g31917,g22003,g31478);
	or 	XG16623 	(g28308,g15795,g27105);
	or 	XG16624 	(g28681,g16634,g27428);
	or 	XG16625 	(g30414,g21794,g30002);
	or 	XG16626 	(g31883,g21777,g31132);
	or 	XG16627 	(g28306,g15794,g27104);
	or 	XG16628 	(g31925,g22061,g31789);
	or 	XG16629 	(g31304,g29608,g29594);
	or 	XG16630 	(g28716,g13887,g27481);
	or 	XG16631 	(g28850,g16869,g27557);
	or 	XG16632 	(g28668,g16617,g27411);
	or 	XG16633 	(g31920,g22045,g31493);
	or 	XG16634 	(g31921,g22046,g31508);
	or 	XG16635 	(g31884,g21778,g31290);
	and 	XG16636 	(g28556,g20374,g27431);
	and 	XG16637 	(g28530,g20240,g27383);
	and 	XG16638 	(g33332,g20608,g32217);
	and 	XG16639 	(g33338,g20633,g32220);
	and 	XG16640 	(g33342,g20660,g32226);
	and 	XG16641 	(g33327,g20561,g32208);
	and 	XG16642 	(g33328,g20584,g32209);
	and 	XG16643 	(g33349,g20699,g32233);
	and 	XG16644 	(g28239,g19659,g27135);
	and 	XG16645 	(g33331,g20607,g32216);
	and 	XG16646 	(g33350,g20702,g32235);
	and 	XG16647 	(g33355,g20769,g32243);
	and 	XG16648 	(g33329,g20585,g32210);
	and 	XG16649 	(g33369,g21060,g32277);
	and 	XG16650 	(g33352,g20712,g32237);
	and 	XG16651 	(g33372,g21183,g32285);
	and 	XG16652 	(g33345,g20671,g32229);
	and 	XG16653 	(g33759,g22847,g33123);
	and 	XG16654 	(g28249,g19677,g27152);
	and 	XG16655 	(g33367,g21053,g32271);
	and 	XG16656 	(g33339,g20634,g32221);
	and 	XG16657 	(g33343,g20665,g32227);
	and 	XG16658 	(g33362,g20914,g32259);
	or 	XG16659 	(g28317,g15805,g27114);
	or 	XG16660 	(g28387,g15858,g27203);
	or 	XG16661 	(g28628,g16531,g27370);
	or 	XG16662 	(g28623,g16520,g27361);
	or 	XG16663 	(g28418,g15882,g27220);
	or 	XG16664 	(g28682,g16635,g27430);
	or 	XG16665 	(g28744,g16759,g27518);
	or 	XG16666 	(g28718,g16702,g27483);
	or 	XG16667 	(g28622,g16519,g27360);
	or 	XG16668 	(g28345,g15821,g27137);
	or 	XG16669 	(g28688,g16639,g27435);
	or 	XG16670 	(g28745,g16760,g27519);
	or 	XG16671 	(g28310,g15797,g27107);
	or 	XG16672 	(g28774,g16804,g27536);
	or 	XG16673 	(g28374,g15850,g27181);
	or 	XG16674 	(g28309,g15796,g27106);
	or 	XG16675 	(g28319,g15807,g27115);
	and 	XG16676 	(g31526,g29342,g22521);
	nand 	XG16677 	(I26440,I26438,g14271);
	or 	XG16678 	(g31259,g29554,g25992);
	or 	XG16679 	(g28729,g16732,g27502);
	or 	XG16680 	(g28430,g15914,g27229);
	or 	XG16681 	(g28636,g16538,g27376);
	or 	XG16682 	(g28772,g16802,g27534);
	or 	XG16683 	(g28667,g16616,g27410);
	or 	XG16684 	(g29143,g17146,g27650);
	or 	XG16685 	(g31260,g29555,g25993);
	or 	XG16686 	(g28773,g16803,g27535);
	or 	XG16687 	(g28701,g16669,g27455);
	or 	XG16688 	(g28296,g15784,g27095);
	or 	XG16689 	(g28746,g16762,g27520);
	or 	XG16690 	(g28511,g16208,g27272);
	or 	XG16691 	(g28429,g15913,g27228);
	or 	XG16692 	(g28719,g16703,g27485);
	or 	XG16693 	(g28708,g16674,g27462);
	or 	XG16694 	(g31251,g29527,g25973);
	or 	XG16695 	(g28749,g16764,g27523);
	or 	XG16696 	(g28730,g13912,g27503);
	or 	XG16697 	(g28419,g15884,g27221);
	or 	XG16698 	(g28700,g16668,g27454);
	or 	XG16699 	(g28732,g16734,g27505);
	or 	XG16700 	(g28389,g15860,g27206);
	or 	XG16701 	(g28671,g16619,g27413);
	or 	XG16702 	(g31772,g28654,g30035);
	or 	XG16703 	(g28751,g16766,g27526);
	or 	XG16704 	(g31322,g29635,g26128);
	or 	XG16705 	(g28643,g16592,g27386);
	or 	XG16706 	(g28634,g16536,g27374);
	not 	XG16707 	(g32186,I29720);
	or 	XG16708 	(g28405,g15875,g27216);
	or 	XG16709 	(g28851,g16870,g27558);
	or 	XG16710 	(g28735,g16737,g27510);
	or 	XG16711 	(g28631,g16534,g27372);
	or 	XG16712 	(g28322,g15809,g27117);
	or 	XG16713 	(g28704,g16671,g27459);
	or 	XG16714 	(g28748,g16763,g27522);
	or 	XG16715 	(g28699,g16667,g27452);
	nand 	XG16716 	(I26072,I26070,g13517);
	or 	XG16717 	(g28817,g16845,g27548);
	or 	XG16718 	(g28724,g16707,g27491);
	or 	XG16719 	(g31473,g29666,g26180);
	or 	XG16720 	(g28687,g16638,g27434);
	or 	XG16721 	(g28690,g16641,g27436);
	nand 	XG16722 	(g34174,g12323,g33851,g617);
	and 	XG16723 	(g34084,g33851,g9214);
	or 	XG16724 	(g31256,g29537,g25983);
	not 	XG16725 	(g34161,g33851);
	nand 	XG16726 	(I26368,I26366,g14211);
	nand 	XG16727 	(I26051,I26049,g13500);
	or 	XG16728 	(g31246,g29518,g25965);
	or 	XG16729 	(g28661,g16611,g27406);
	or 	XG16730 	(g28650,g16598,g27391);
	or 	XG16731 	(g28670,g16618,g27412);
	or 	XG16732 	(g28818,g13998,g27549);
	or 	XG16733 	(g28884,g16885,g27568);
	or 	XG16734 	(g28777,g16807,g27539);
	nand 	XG16735 	(I26095,I26093,g13539);
	or 	XG16736 	(g31466,g29650,g26160);
	or 	XG16737 	(g31250,g29526,g25972);
	or 	XG16738 	(g33964,g18146,g33817);
	or 	XG16739 	(g33542,g18265,g33102);
	and 	XG16740 	(g34071,g33799,g8854);
	or 	XG16741 	(g33534,g21700,g33186);
	or 	XG16742 	(g33536,g21715,g33241);
	or 	XG16743 	(g33539,g18178,g33245);
	or 	XG16744 	(g33540,g18207,g33099);
	or 	XG16745 	(g34125,g33124,g33724);
	or 	XG16746 	(g33788,g32041,g33122);
	and 	XG16747 	(g28588,g20499,g27489);
	and 	XG16748 	(g33873,g20549,g33291);
	and 	XG16749 	(g33356,g20772,g32245);
	and 	XG16750 	(g33361,g20911,g32257);
	and 	XG16751 	(g34157,g20159,g33794);
	and 	XG16752 	(g33805,g20079,g33232);
	and 	XG16753 	(g28252,g19682,g27159);
	and 	XG16754 	(g28571,g20435,g27458);
	or 	XG16755 	(g33535,g21711,g33233);
	or 	XG16756 	(g33537,g21716,g33244);
	or 	XG16757 	(g33732,g32011,g33104);
	not 	XG16758 	(g33797,g33306);
	nor 	XG16759 	(g33823,g11083,g33306,g8774);
	and 	XG16760 	(g33717,g33306,g14092);
	and 	XG16761 	(g33710,g33246,g14037);
	and 	XG16762 	(g33789,g23022,g33159);
	or 	XG16763 	(g33608,g18537,g33322);
	or 	XG16764 	(g33733,g32012,g33105);
	nor 	XG16765 	(g30601,g29718,g16279);
	or 	XG16766 	(g30672,g29752,g13737);
	not 	XG16767 	(g30237,I28480);
	not 	XG16768 	(g30259,g28463);
	not 	XG16769 	(g30206,g28436);
	and 	XG16770 	(g31994,g22215,g31775);
	and 	XG16771 	(g31989,g22200,g31770);
	and 	XG16772 	(g31975,g22177,g31761);
	and 	XG16773 	(g31961,g22154,g31751);
	and 	XG16774 	(g32302,g23485,g31279);
	and 	XG16775 	(g32313,g23515,g31303);
	and 	XG16776 	(g31992,g22213,g31773);
	and 	XG16777 	(g31505,g24379,g30195);
	and 	XG16778 	(g31944,g22146,g31745);
	and 	XG16779 	(g32311,g20582,g31295);
	and 	XG16780 	(g32232,g20266,g31241);
	and 	XG16781 	(g32281,g20500,g31257);
	and 	XG16782 	(g32325,g23538,g31316);
	and 	XG16783 	(g32255,g20381,g31248);
	and 	XG16784 	(g32290,g20525,g31267);
	and 	XG16785 	(g32008,g22223,g31781);
	and 	XG16786 	(g32340,g23585,g31468);
	and 	XG16787 	(g32337,g20663,g31465);
	and 	XG16788 	(g32270,g20444,g31254);
	and 	XG16789 	(g32282,g20503,g31258);
	or 	XG16790 	(I30261,g30825,g30735,g31376,g29385);
	or 	XG16791 	(I30192,g30825,g30735,g31376,g29385);
	or 	XG16792 	(I29985,g30825,g30735,g31376,g29385);
	or 	XG16793 	(I30123,g30825,g30735,g31376,g29385);
	or 	XG16794 	(I30468,g30825,g30735,g31376,g29385);
	or 	XG16795 	(I30054,g30825,g30735,g31376,g29385);
	or 	XG16796 	(I30399,g30825,g30735,g31376,g29385);
	or 	XG16797 	(I30330,g30825,g30735,g31376,g29385);
	not 	XG16798 	(g32118,g31008);
	not 	XG16799 	(g32033,g30929);
	not 	XG16800 	(g32038,g30934);
	or 	XG16801 	(g33259,g29521,g32109);
	and 	XG16802 	(g32030,g30937,g4172);
	or 	XG16803 	(g33251,g29509,g32096);
	and 	XG16804 	(g32303,g31376,g27550);
	or 	XG16805 	(g30609,g29742,g13633);
	and 	XG16806 	(g32335,g31566,g6199);
	not 	XG16807 	(g28954,g27830);
	and 	XG16808 	(g32328,g31554,g5853);
	and 	XG16809 	(g32410,g30997,g4933);
	and 	XG16810 	(g32317,g31542,g5507);
	not 	XG16811 	(I26700,g27956);
	and 	XG16812 	(g31933,g30735,g939);
	not 	XG16813 	(I26693,g27930);
	and 	XG16814 	(g32069,g30735,g10878);
	not 	XG16815 	(I27481,g27928);
	and 	XG16816 	(g32167,g31194,g3853);
	and 	XG16817 	(g31985,g30614,g4722);
	or 	XG16818 	(g33279,g29573,g32140);
	and 	XG16819 	(g32013,g30614,g8673);
	and 	XG16820 	(g32309,g31528,g5160);
	and 	XG16821 	(g32095,g30825,g7619);
	and 	XG16822 	(g32161,g31154,g3151);
	and 	XG16823 	(g32409,g30996,g4754);
	and 	XG16824 	(g32047,g31070,g27248);
	or 	XG16825 	(g30734,g29774,g13808);
	or 	XG16826 	(g32266,g29354,g30604);
	and 	XG16827 	(g32014,g30673,g8715);
	and 	XG16828 	(g32088,g31070,g27241);
	and 	XG16829 	(g32056,g31021,g27271);
	or 	XG16830 	(g33380,g29926,g32234);
	or 	XG16831 	(g30608,g29736,g13604);
	and 	XG16832 	(g32082,g30673,g4917);
	and 	XG16833 	(g32054,g30735,g10890);
	not 	XG16834 	(g31771,I29337);
	and 	XG16835 	(g32402,g30990,g4888);
	and 	XG16836 	(g31941,g30825,g1283);
	or 	XG16837 	(g30611,g29743,g13671);
	or 	XG16838 	(I30193,g31528,g30673,g30614,g31070);
	or 	XG16839 	(I30055,g30673,g30614,g31170,g31070);
	or 	XG16840 	(I29986,g30673,g30614,g31194,g31070);
	or 	XG16841 	(I30124,g30673,g30614,g31154,g31070);
	not 	XG16842 	(g32462,g30673);
	not 	XG16843 	(g32534,g30673);
	not 	XG16844 	(g32649,g30673);
	not 	XG16845 	(g32541,g30673);
	not 	XG16846 	(g32613,g30673);
	not 	XG16847 	(g32584,g30673);
	not 	XG16848 	(g32519,g30673);
	not 	XG16849 	(g32555,g30673);
	not 	XG16850 	(g32476,g30673);
	not 	XG16851 	(g32874,g30673);
	not 	XG16852 	(g32853,g30673);
	not 	XG16853 	(g32713,g30673);
	not 	XG16854 	(g32656,g30673);
	not 	XG16855 	(g32599,g30673);
	not 	XG16856 	(g32504,g30673);
	not 	XG16857 	(g32548,g30673);
	not 	XG16858 	(g32627,g30673);
	not 	XG16859 	(g32620,g30673);
	not 	XG16860 	(g32881,g30673);
	not 	XG16861 	(g32691,g30673);
	not 	XG16862 	(g32592,g30673);
	not 	XG16863 	(g32634,g30673);
	not 	XG16864 	(g32483,g30673);
	not 	XG16865 	(g32663,g30673);
	not 	XG16866 	(g32606,g30673);
	not 	XG16867 	(g32684,g30673);
	not 	XG16868 	(g32569,g30673);
	not 	XG16869 	(g32677,g30673);
	not 	XG16870 	(g32469,g30673);
	not 	XG16871 	(g32670,g30673);
	not 	XG16872 	(g32706,g30673);
	not 	XG16873 	(g32867,g30673);
	not 	XG16874 	(g32527,g30673);
	not 	XG16875 	(g32497,g30673);
	not 	XG16876 	(g32860,g30673);
	not 	XG16877 	(g32888,g30673);
	not 	XG16878 	(g32490,g30673);
	not 	XG16879 	(g32895,g30673);
	not 	XG16880 	(g32562,g30673);
	not 	XG16881 	(g32902,g30673);
	not 	XG16882 	(g32754,g30825);
	not 	XG16883 	(g32472,g30825);
	not 	XG16884 	(g32573,g30825);
	not 	XG16885 	(g32718,g30825);
	not 	XG16886 	(g32898,g30825);
	not 	XG16887 	(g32927,g30825);
	not 	XG16888 	(g32682,g30825);
	not 	XG16889 	(g32920,g30825);
	not 	XG16890 	(g32812,g30825);
	not 	XG16891 	(g32833,g30825);
	not 	XG16892 	(g32848,g30825);
	not 	XG16893 	(g32725,g30825);
	not 	XG16894 	(g32515,g30825);
	not 	XG16895 	(g32761,g30825);
	not 	XG16896 	(g32732,g30825);
	not 	XG16897 	(g32963,g30825);
	not 	XG16898 	(g32653,g30825);
	not 	XG16899 	(g32566,g30825);
	not 	XG16900 	(g32501,g30825);
	not 	XG16901 	(g32588,g30825);
	not 	XG16902 	(g32494,g30825);
	not 	XG16903 	(g32595,g30825);
	not 	XG16904 	(g32617,g30825);
	not 	XG16905 	(g32559,g30825);
	not 	XG16906 	(g32631,g30825);
	not 	XG16907 	(g32783,g30825);
	not 	XG16908 	(g32458,g30825);
	not 	XG16909 	(g32970,g30825);
	not 	XG16910 	(g32602,g30825);
	not 	XG16911 	(g32696,g30825);
	not 	XG16912 	(g32775,g30825);
	not 	XG16913 	(g32826,g30825);
	not 	XG16914 	(g32552,g30825);
	not 	XG16915 	(g32710,g30825);
	not 	XG16916 	(g32768,g30825);
	not 	XG16917 	(g32508,g30825);
	not 	XG16918 	(g32949,g30825);
	not 	XG16919 	(g32862,g30825);
	not 	XG16920 	(g32840,g30825);
	not 	XG16921 	(g32537,g30825);
	not 	XG16922 	(g32891,g30825);
	not 	XG16923 	(g32797,g30825);
	not 	XG16924 	(g32530,g30825);
	not 	XG16925 	(g32905,g30825);
	not 	XG16926 	(g32913,g30825);
	not 	XG16927 	(g32790,g30825);
	not 	XG16928 	(g32703,g30825);
	not 	XG16929 	(g32523,g30825);
	not 	XG16930 	(g32465,g30825);
	not 	XG16931 	(g32638,g30825);
	not 	XG16932 	(g32747,g30825);
	not 	XG16933 	(g32580,g30825);
	not 	XG16934 	(g32884,g30825);
	not 	XG16935 	(g32487,g30825);
	not 	XG16936 	(g32667,g30825);
	not 	XG16937 	(g32942,g30825);
	not 	XG16938 	(g32660,g30825);
	not 	XG16939 	(g32624,g30825);
	not 	XG16940 	(g32689,g30825);
	not 	XG16941 	(g32877,g30825);
	not 	XG16942 	(g32819,g30825);
	not 	XG16943 	(g32855,g30825);
	not 	XG16944 	(g32956,g30825);
	not 	XG16945 	(g32645,g30825);
	or 	XG16946 	(I30400,g30614,g31327,g30937,g31021);
	not 	XG16947 	(g32859,g30614);
	not 	XG16948 	(g32591,g30614);
	not 	XG16949 	(g32612,g30614);
	not 	XG16950 	(g32648,g30614);
	not 	XG16951 	(g32605,g30614);
	not 	XG16952 	(g32683,g30614);
	not 	XG16953 	(g32554,g30614);
	not 	XG16954 	(g32576,g30614);
	not 	XG16955 	(g32852,g30614);
	not 	XG16956 	(g32518,g30614);
	not 	XG16957 	(g32712,g30614);
	not 	XG16958 	(g32705,g30614);
	not 	XG16959 	(g32489,g30614);
	not 	XG16960 	(g32669,g30614);
	not 	XG16961 	(g32561,g30614);
	not 	XG16962 	(g32598,g30614);
	not 	XG16963 	(g32887,g30614);
	not 	XG16964 	(g32461,g30614);
	not 	XG16965 	(g32880,g30614);
	not 	XG16966 	(g32533,g30614);
	not 	XG16967 	(g32626,g30614);
	not 	XG16968 	(g32482,g30614);
	not 	XG16969 	(g32662,g30614);
	not 	XG16970 	(g32583,g30614);
	not 	XG16971 	(g32641,g30614);
	not 	XG16972 	(g32873,g30614);
	not 	XG16973 	(g32475,g30614);
	not 	XG16974 	(g32909,g30614);
	not 	XG16975 	(g32676,g30614);
	not 	XG16976 	(g32468,g30614);
	not 	XG16977 	(g32619,g30614);
	not 	XG16978 	(g32655,g30614);
	not 	XG16979 	(g32511,g30614);
	not 	XG16980 	(g32866,g30614);
	not 	XG16981 	(g32526,g30614);
	not 	XG16982 	(g32496,g30614);
	not 	XG16983 	(g32894,g30614);
	not 	XG16984 	(g32547,g30614);
	not 	XG16985 	(g32698,g30614);
	not 	XG16986 	(g32540,g30614);
	not 	XG16987 	(I26682,g27774);
	and 	XG16988 	(g32071,g31070,g27236);
	or 	XG16989 	(g30733,g29773,g13807);
	and 	XG16990 	(g32097,g31021,g25960);
	and 	XG16991 	(g32348,g31672,g2145);
	not 	XG16992 	(g29042,I27388);
	and 	XG16993 	(g32086,g30735,g7597);
	not 	XG16994 	(g29372,I27738);
	not 	XG16995 	(I26705,g27967);
	not 	XG16996 	(g28752,I27232);
	and 	XG16997 	(g32342,g31579,g6545);
	and 	XG16998 	(g32369,g31672,g2130);
	not 	XG16999 	(g32858,g31327);
	not 	XG17000 	(g32946,g31327);
	not 	XG17001 	(g32788,g31327);
	not 	XG17002 	(g32795,g31327);
	not 	XG17003 	(g32744,g31327);
	not 	XG17004 	(g32758,g31327);
	not 	XG17005 	(g32809,g31327);
	not 	XG17006 	(g32837,g31327);
	not 	XG17007 	(g32939,g31327);
	not 	XG17008 	(g32865,g31327);
	not 	XG17009 	(g32830,g31327);
	not 	XG17010 	(g32816,g31327);
	not 	XG17011 	(g32823,g31327);
	not 	XG17012 	(g32901,g31327);
	not 	XG17013 	(g32918,g31327);
	not 	XG17014 	(g32967,g31327);
	not 	XG17015 	(g32886,g31327);
	not 	XG17016 	(g32879,g31327);
	not 	XG17017 	(g32960,g31327);
	not 	XG17018 	(g32737,g31327);
	not 	XG17019 	(g32765,g31327);
	not 	XG17020 	(g32730,g31327);
	not 	XG17021 	(g32802,g31327);
	not 	XG17022 	(g32925,g31327);
	not 	XG17023 	(g32723,g31327);
	not 	XG17024 	(g32932,g31327);
	not 	XG17025 	(g32872,g31327);
	not 	XG17026 	(g32851,g31327);
	not 	XG17027 	(g32772,g31327);
	not 	XG17028 	(g32751,g31327);
	not 	XG17029 	(g32908,g31327);
	not 	XG17030 	(g32953,g31327);
	not 	XG17031 	(g32633,g31154);
	not 	XG17032 	(g32604,g31154);
	not 	XG17033 	(g32611,g31154);
	not 	XG17034 	(g32647,g31154);
	not 	XG17035 	(g32640,g31154);
	not 	XG17036 	(g32618,g31154);
	not 	XG17037 	(g32597,g31154);
	not 	XG17038 	(g32590,g31154);
	not 	XG17039 	(g32467,g31194);
	not 	XG17040 	(g32460,g31194);
	not 	XG17041 	(g32488,g31194);
	not 	XG17042 	(g32474,g31194);
	not 	XG17043 	(g32517,g31194);
	not 	XG17044 	(g32510,g31194);
	not 	XG17045 	(g32503,g31194);
	not 	XG17046 	(g32481,g31194);
	not 	XG17047 	(g32539,g31170);
	not 	XG17048 	(g32525,g31170);
	not 	XG17049 	(g32532,g31170);
	not 	XG17050 	(g32582,g31170);
	not 	XG17051 	(g32553,g31170);
	not 	XG17052 	(g32575,g31170);
	not 	XG17053 	(g32568,g31170);
	not 	XG17054 	(g32546,g31170);
	or 	XG17055 	(I30331,g30937,g31021,g31710,g31672);
	or 	XG17056 	(I30469,g30937,g31021,g31710,g31672);
	or 	XG17057 	(I30262,g30937,g31021,g31710,g31672);
	not 	XG17058 	(g32785,g31710);
	not 	XG17059 	(g32777,g31710);
	not 	XG17060 	(g32770,g31710);
	not 	XG17061 	(g32828,g31710);
	not 	XG17062 	(g32972,g31710);
	not 	XG17063 	(g32813,g31710);
	not 	XG17064 	(g32799,g31710);
	not 	XG17065 	(g32748,g31710);
	not 	XG17066 	(g32915,g31710);
	not 	XG17067 	(g32842,g31710);
	not 	XG17068 	(g32792,g31710);
	not 	XG17069 	(g32958,g31710);
	not 	XG17070 	(g32929,g31710);
	not 	XG17071 	(g32727,g31710);
	not 	XG17072 	(g32806,g31710);
	not 	XG17073 	(g32720,g31710);
	not 	XG17074 	(g32835,g31710);
	not 	XG17075 	(g32936,g31710);
	not 	XG17076 	(g32922,g31710);
	not 	XG17077 	(g32965,g31710);
	not 	XG17078 	(g32734,g31710);
	not 	XG17079 	(g32763,g31710);
	not 	XG17080 	(g32741,g31710);
	not 	XG17081 	(g32943,g31710);
	not 	XG17082 	(g32665,g31579);
	not 	XG17083 	(g32693,g31579);
	not 	XG17084 	(g32686,g31579);
	not 	XG17085 	(g32679,g31579);
	not 	XG17086 	(g32672,g31579);
	not 	XG17087 	(g32707,g31579);
	not 	XG17088 	(g32658,g31579);
	not 	XG17089 	(g32700,g31579);
	not 	XG17090 	(g32628,g31542);
	not 	XG17091 	(g32642,g31542);
	not 	XG17092 	(g32621,g31542);
	not 	XG17093 	(g32635,g31542);
	not 	XG17094 	(g32593,g31542);
	not 	XG17095 	(g32607,g31542);
	not 	XG17096 	(g32614,g31542);
	not 	XG17097 	(g32600,g31542);
	not 	XG17098 	(g32950,g31672);
	not 	XG17099 	(g32776,g31672);
	not 	XG17100 	(g32719,g31672);
	not 	XG17101 	(g32755,g31672);
	not 	XG17102 	(g32805,g31672);
	not 	XG17103 	(g32798,g31672);
	not 	XG17104 	(g32921,g31672);
	not 	XG17105 	(g32935,g31672);
	not 	XG17106 	(g32914,g31672);
	not 	XG17107 	(g32733,g31672);
	not 	XG17108 	(g32971,g31672);
	not 	XG17109 	(g32769,g31672);
	not 	XG17110 	(g32827,g31672);
	not 	XG17111 	(g32928,g31672);
	not 	XG17112 	(g32820,g31672);
	not 	XG17113 	(g32726,g31672);
	not 	XG17114 	(g32834,g31672);
	not 	XG17115 	(g32841,g31672);
	not 	XG17116 	(g32964,g31672);
	not 	XG17117 	(g32762,g31672);
	not 	XG17118 	(g32740,g31672);
	not 	XG17119 	(g32791,g31672);
	not 	XG17120 	(g32784,g31672);
	not 	XG17121 	(g32957,g31672);
	not 	XG17122 	(g32692,g31528);
	not 	XG17123 	(g32664,g31528);
	not 	XG17124 	(g32678,g31528);
	not 	XG17125 	(g32657,g31528);
	not 	XG17126 	(g32685,g31528);
	not 	XG17127 	(g32714,g31528);
	not 	XG17128 	(g32671,g31528);
	not 	XG17129 	(g32699,g31528);
	not 	XG17130 	(g32491,g31566);
	not 	XG17131 	(g32463,g31566);
	not 	XG17132 	(g32484,g31566);
	not 	XG17133 	(g32477,g31566);
	not 	XG17134 	(g32470,g31566);
	not 	XG17135 	(g32498,g31566);
	not 	XG17136 	(g32512,g31566);
	not 	XG17137 	(g32505,g31566);
	not 	XG17138 	(g32563,g31554);
	not 	XG17139 	(g32535,g31554);
	not 	XG17140 	(g32577,g31554);
	not 	XG17141 	(g32570,g31554);
	not 	XG17142 	(g32528,g31554);
	not 	XG17143 	(g32549,g31554);
	not 	XG17144 	(g32542,g31554);
	not 	XG17145 	(g32556,g31554);
	not 	XG17146 	(g32899,g31021);
	not 	XG17147 	(g32951,g31021);
	not 	XG17148 	(g32849,g31021);
	not 	XG17149 	(g32771,g31021);
	not 	XG17150 	(g32973,g31021);
	not 	XG17151 	(g32906,g31021);
	not 	XG17152 	(g32728,g31021);
	not 	XG17153 	(g32892,g31021);
	not 	XG17154 	(g32749,g31021);
	not 	XG17155 	(g32836,g31021);
	not 	XG17156 	(g32966,g31021);
	not 	XG17157 	(g32843,g31021);
	not 	XG17158 	(g32856,g31021);
	not 	XG17159 	(g32793,g31021);
	not 	XG17160 	(g32944,g31021);
	not 	XG17161 	(g32742,g31021);
	not 	XG17162 	(g32786,g31021);
	not 	XG17163 	(g32778,g31021);
	not 	XG17164 	(g32756,g31021);
	not 	XG17165 	(g32821,g31021);
	not 	XG17166 	(g32863,g31021);
	not 	XG17167 	(g32807,g31021);
	not 	XG17168 	(g32814,g31021);
	not 	XG17169 	(g32800,g31021);
	not 	XG17170 	(g32937,g31021);
	not 	XG17171 	(g32930,g31021);
	not 	XG17172 	(g32721,g31021);
	not 	XG17173 	(g32916,g31021);
	not 	XG17174 	(g32885,g31021);
	not 	XG17175 	(g32923,g31021);
	not 	XG17176 	(g32735,g31021);
	not 	XG17177 	(g32870,g31021);
	not 	XG17178 	(g32844,g30937);
	not 	XG17179 	(g32871,g30937);
	not 	XG17180 	(g32794,g30937);
	not 	XG17181 	(g32829,g30937);
	not 	XG17182 	(g32729,g30937);
	not 	XG17183 	(g32907,g30937);
	not 	XG17184 	(g32808,g30937);
	not 	XG17185 	(g32900,g30937);
	not 	XG17186 	(g32864,g30937);
	not 	XG17187 	(g32822,g30937);
	not 	XG17188 	(g32938,g30937);
	not 	XG17189 	(g32893,g30937);
	not 	XG17190 	(g32878,g30937);
	not 	XG17191 	(g32764,g30937);
	not 	XG17192 	(g32736,g30937);
	not 	XG17193 	(g32924,g30937);
	not 	XG17194 	(g32722,g30937);
	not 	XG17195 	(g32857,g30937);
	not 	XG17196 	(g32959,g30937);
	not 	XG17197 	(g32850,g30937);
	not 	XG17198 	(g32945,g30937);
	not 	XG17199 	(g32779,g30937);
	not 	XG17200 	(g32743,g30937);
	not 	XG17201 	(g32787,g30937);
	not 	XG17202 	(g32757,g30937);
	not 	XG17203 	(g32750,g30937);
	not 	XG17204 	(g32952,g30937);
	not 	XG17205 	(g32974,g30937);
	not 	XG17206 	(g32815,g30937);
	not 	XG17207 	(g32917,g30937);
	not 	XG17208 	(g32801,g30937);
	not 	XG17209 	(g32931,g30937);
	not 	XG17210 	(g32473,g31070);
	not 	XG17211 	(g32538,g31070);
	not 	XG17212 	(g32675,g31070);
	not 	XG17213 	(g32567,g31070);
	not 	XG17214 	(g32560,g31070);
	not 	XG17215 	(g32466,g31070);
	not 	XG17216 	(g32704,g31070);
	not 	XG17217 	(g32524,g31070);
	not 	XG17218 	(g32589,g31070);
	not 	XG17219 	(g32610,g31070);
	not 	XG17220 	(g32668,g31070);
	not 	XG17221 	(g32495,g31070);
	not 	XG17222 	(g32545,g31070);
	not 	XG17223 	(g32459,g31070);
	not 	XG17224 	(g32697,g31070);
	not 	XG17225 	(g32690,g31070);
	not 	XG17226 	(g32603,g31070);
	not 	XG17227 	(g32646,g31070);
	not 	XG17228 	(g32574,g31070);
	not 	XG17229 	(g32509,g31070);
	not 	XG17230 	(g32711,g31070);
	not 	XG17231 	(g32516,g31070);
	not 	XG17232 	(g32639,g31070);
	not 	XG17233 	(g32654,g31070);
	not 	XG17234 	(g32531,g31070);
	not 	XG17235 	(g32502,g31070);
	not 	XG17236 	(g32596,g31070);
	not 	XG17237 	(g32480,g31070);
	not 	XG17238 	(g32581,g31070);
	not 	XG17239 	(g32625,g31070);
	not 	XG17240 	(g32661,g31070);
	not 	XG17241 	(g32632,g31070);
	or 	XG17242 	(g33255,g29514,g32106);
	or 	XG17243 	(g32251,g29352,g30599);
	not 	XG17244 	(g28779,I27253);
	and 	XG17245 	(g32321,g31376,g27613);
	and 	XG17246 	(g32400,g30989,g4743);
	or 	XG17247 	(g30605,g29520,g29529);
	or 	XG17248 	(g30597,g29693,g13564);
	nand 	XG17249 	(g32057,g13297,g31003);
	not 	XG17250 	(I26676,g27736);
	and 	XG17251 	(g32414,g30999,g4944);
	or 	XG17252 	(g33274,g29563,g32126);
	not 	XG17253 	(I28585,g30217);
	or 	XG17254 	(g29539,g28220,g2864);
	or 	XG17255 	(g32231,g29346,g30590);
	and 	XG17256 	(g32295,g31376,g27931);
	and 	XG17257 	(I31593,g7788,g8350,g31003);
	not 	XG17258 	(g32099,g31009);
	not 	XG17259 	(g32090,g31003);
	not 	XG17260 	(I27271,g27998);
	not 	XG17261 	(g30591,I28851);
	or 	XG17262 	(I28147,g28220,g24561,g2946);
	not 	XG17263 	(g28917,I27314);
	not 	XG17264 	(I27784,g29013);
	and 	XG17265 	(g32200,g31376,g27468);
	not 	XG17266 	(I26785,g27013);
	and 	XG17267 	(g32196,g31376,g27587);
	or 	XG17268 	(g30317,I28567,I28566,g29208);
	not 	XG17269 	(g28367,I26880);
	not 	XG17270 	(I26670,g27709);
	not 	XG17271 	(I27777,g29043);
	not 	XG17272 	(I26679,g27773);
	and 	XG17273 	(g32049,g30735,g10902);
	not 	XG17274 	(I26687,g27880);
	not 	XG17275 	(I26649,g27675);
	not 	XG17276 	(I28419,g29195);
	and 	XG17277 	(g32046,g30735,g10925);
	and 	XG17278 	(g32191,g31376,g27593);
	or 	XG17279 	(g32239,g29350,g30595);
	not 	XG17280 	(g32825,g30735);
	not 	XG17281 	(g32832,g30735);
	not 	XG17282 	(g32767,g30735);
	not 	XG17283 	(g32760,g30735);
	not 	XG17284 	(g32724,g30735);
	not 	XG17285 	(g32789,g30735);
	not 	XG17286 	(g32507,g30735);
	not 	XG17287 	(g32514,g30735);
	not 	XG17288 	(g32500,g30735);
	not 	XG17289 	(g32962,g30735);
	not 	XG17290 	(g32804,g30735);
	not 	XG17291 	(g32652,g30735);
	not 	XG17292 	(g32934,g30735);
	not 	XG17293 	(g32674,g30735);
	not 	XG17294 	(g32609,g30735);
	not 	XG17295 	(g32883,g30735);
	not 	XG17296 	(g32637,g30735);
	not 	XG17297 	(g32941,g30735);
	not 	XG17298 	(g32594,g30735);
	not 	XG17299 	(g32630,g30735);
	not 	XG17300 	(g32616,g30735);
	not 	XG17301 	(g32782,g30735);
	not 	XG17302 	(g32623,g30735);
	not 	XG17303 	(g32544,g30735);
	not 	XG17304 	(g32558,g30735);
	not 	XG17305 	(g32919,g30735);
	not 	XG17306 	(g32955,g30735);
	not 	XG17307 	(g32774,g30735);
	not 	XG17308 	(g32709,g30735);
	not 	XG17309 	(g32869,g30735);
	not 	XG17310 	(g32529,g30735);
	not 	XG17311 	(g32753,g30735);
	not 	XG17312 	(g32681,g30735);
	not 	XG17313 	(g32811,g30735);
	not 	XG17314 	(g32717,g30735);
	not 	XG17315 	(g32897,g30735);
	not 	XG17316 	(g32890,g30735);
	not 	XG17317 	(g32912,g30735);
	not 	XG17318 	(g32847,g30735);
	not 	XG17319 	(g32904,g30735);
	not 	XG17320 	(g32702,g30735);
	not 	XG17321 	(g32948,g30735);
	not 	XG17322 	(g32522,g30735);
	not 	XG17323 	(g32464,g30735);
	not 	XG17324 	(g32565,g30735);
	not 	XG17325 	(g32493,g30735);
	not 	XG17326 	(g32746,g30735);
	not 	XG17327 	(g32579,g30735);
	not 	XG17328 	(g32587,g30735);
	not 	XG17329 	(g32486,g30735);
	not 	XG17330 	(g32479,g30735);
	not 	XG17331 	(g32839,g30735);
	not 	XG17332 	(g32854,g30735);
	not 	XG17333 	(g32876,g30735);
	not 	XG17334 	(g32688,g30735);
	not 	XG17335 	(g32457,g30735);
	not 	XG17336 	(g32695,g30735);
	not 	XG17337 	(g32818,g30735);
	not 	XG17338 	(g32969,g30735);
	not 	XG17339 	(g32644,g30735);
	not 	XG17340 	(g32659,g30735);
	not 	XG17341 	(g32572,g30735);
	not 	XG17342 	(g32551,g30735);
	not 	XG17343 	(g32739,g30735);
	not 	XG17344 	(g32911,g31376);
	not 	XG17345 	(g32629,g31376);
	not 	XG17346 	(g32766,g31376);
	not 	XG17347 	(g32701,g31376);
	not 	XG17348 	(g32926,g31376);
	not 	XG17349 	(g32861,g31376);
	not 	XG17350 	(g32521,g31376);
	not 	XG17351 	(g32903,g31376);
	not 	XG17352 	(g32506,g31376);
	not 	XG17353 	(g32947,g31376);
	not 	XG17354 	(g32940,g31376);
	not 	XG17355 	(g32759,g31376);
	not 	XG17356 	(g32882,g31376);
	not 	XG17357 	(g32745,g31376);
	not 	XG17358 	(g32608,g31376);
	not 	XG17359 	(g32636,g31376);
	not 	XG17360 	(g32622,g31376);
	not 	XG17361 	(g32485,g31376);
	not 	XG17362 	(g32875,g31376);
	not 	XG17363 	(g32643,g31376);
	not 	XG17364 	(g32954,g31376);
	not 	XG17365 	(g32752,g31376);
	not 	XG17366 	(g32687,g31376);
	not 	XG17367 	(g32571,g31376);
	not 	XG17368 	(g32680,g31376);
	not 	XG17369 	(g32817,g31376);
	not 	XG17370 	(g32810,g31376);
	not 	XG17371 	(g32471,g31376);
	not 	XG17372 	(g32708,g31376);
	not 	XG17373 	(g32868,g31376);
	not 	XG17374 	(g32499,g31376);
	not 	XG17375 	(g32831,g31376);
	not 	XG17376 	(g32716,g31376);
	not 	XG17377 	(g32896,g31376);
	not 	XG17378 	(g32961,g31376);
	not 	XG17379 	(g32513,g31376);
	not 	XG17380 	(g32651,g31376);
	not 	XG17381 	(g32803,g31376);
	not 	XG17382 	(g32731,g31376);
	not 	XG17383 	(g32846,g31376);
	not 	XG17384 	(g32933,g31376);
	not 	XG17385 	(g32673,g31376);
	not 	XG17386 	(g32564,g31376);
	not 	XG17387 	(g32536,g31376);
	not 	XG17388 	(g32796,g31376);
	not 	XG17389 	(g32492,g31376);
	not 	XG17390 	(g32781,g31376);
	not 	XG17391 	(g32615,g31376);
	not 	XG17392 	(g32586,g31376);
	not 	XG17393 	(g32578,g31376);
	not 	XG17394 	(g32543,g31376);
	not 	XG17395 	(g32478,g31376);
	not 	XG17396 	(g32666,g31376);
	not 	XG17397 	(g32601,g31376);
	not 	XG17398 	(g32557,g31376);
	not 	XG17399 	(g32838,g31376);
	not 	XG17400 	(g32694,g31376);
	not 	XG17401 	(g32773,g31376);
	not 	XG17402 	(g32550,g31376);
	not 	XG17403 	(g32456,g31376);
	not 	XG17404 	(g32968,g31376);
	not 	XG17405 	(g32824,g31376);
	not 	XG17406 	(g32889,g31376);
	not 	XG17407 	(g32738,g31376);
	not 	XG17408 	(I26664,g27708);
	not 	XG17409 	(g31596,I29204);
	not 	XG17410 	(I27385,g27438);
	or 	XG17411 	(g33266,g29532,g32114);
	and 	XG17412 	(g32224,g31327,g4300);
	nor 	XG17413 	(g30613,g29365,g4507);
	or 	XG17414 	(g33596,g18494,g33341);
	and 	XG17415 	(g32188,g31376,g27586);
	or 	XG17416 	(g33303,g29638,g32159);
	nor 	XG17417 	(g30922,g29810,g16662);
	nor 	XG17418 	(g29873,g28458,g6875);
	and 	XG17419 	(g32198,g31327,g4253);
	or 	XG17420 	(g30916,g29799,g13853);
	and 	XG17421 	(g32050,g30825,g11003);
	and 	XG17422 	(g32356,g31710,g2704);
	and 	XG17423 	(g31940,g30735,g943);
	and 	XG17424 	(g32396,g30983,g4698);
	nor 	XG17425 	(g30271,g29008,g7041);
	and 	XG17426 	(g30315,g5644,g7028,g29182);
	nor 	XG17427 	(g30262,g29008,g5644);
	and 	XG17428 	(g32350,g31710,g2697);
	or 	XG17429 	(g33597,g18495,g33344);
	or 	XG17430 	(g33383,g29940,g32244);
	and 	XG17431 	(g31502,g29311,g2472);
	and 	XG17432 	(g32310,g31376,g27577);
	nor 	XG17433 	(g30252,g29008,g7028);
	or 	XG17434 	(g33267,g29535,g32115);
	and 	XG17435 	(g32083,g30735,g947);
	or 	XG17436 	(g33254,g29512,g32104);
	and 	XG17437 	(g32176,g31623,g2779);
	not 	XG17438 	(g31522,I29185);
	and 	XG17439 	(g31943,g30614,g4717);
	or 	XG17440 	(g33265,g29530,g32113);
	or 	XG17441 	(g33386,g29951,g32258);
	or 	XG17442 	(g33282,g29577,g32143);
	and 	XG17443 	(g32067,g30614,g4727);
	or 	XG17444 	(g33286,g29585,g32145);
	or 	XG17445 	(g33288,g29587,g32147);
	not 	XG17446 	(g31189,I29002);
	or 	XG17447 	(g33595,g18489,g33368);
	and 	XG17448 	(g32293,g30593,g2827);
	not 	XG17449 	(g31213,I29013);
	or 	XG17450 	(g33277,g29568,g32129);
	or 	XG17451 	(g33384,g29943,g32248);
	and 	XG17452 	(g31480,g30296,g1644);
	and 	XG17453 	(g32376,g31710,g2689);
	and 	XG17454 	(g32204,g31327,g4245);
	and 	XG17455 	(g32172,g31608,g2767);
	nand 	XG17456 	(g32072,g13301,g31009);
	or 	XG17457 	(g33272,g29551,g32121);
	or 	XG17458 	(g33295,g29605,g32153);
	or 	XG17459 	(g30732,g29762,g13778);
	and 	XG17460 	(g31495,g30309,g1913);
	and 	XG17461 	(g32412,g30998,g4765);
	and 	XG17462 	(g32035,g30937,g4176);
	and 	XG17463 	(g32203,g31327,g4249);
	or 	XG17464 	(g33256,g29517,g32107);
	or 	XG17465 	(g33287,g29586,g32146);
	or 	XG17466 	(g33290,g29589,g32149);
	or 	XG17467 	(g33297,g29621,g32157);
	and 	XG17468 	(g32087,g30825,g1291);
	and 	XG17469 	(g32180,g31638,g2791);
	and 	XG17470 	(g31496,g30312,g2338);
	and 	XG17471 	(g32345,g31672,g2138);
	and 	XG17472 	(I31600,g7809,g8400,g31009);
	and 	XG17473 	(g31949,g30825,g1287);
	or 	XG17474 	(g33271,g29549,g32120);
	and 	XG17475 	(g32419,g31000,g4955);
	or 	XG17476 	(g33581,g18443,g33333);
	or 	XG17477 	(g33298,g29622,g32158);
	or 	XG17478 	(g33273,g29553,g32122);
	or 	XG17479 	(g33278,g29572,g32139);
	and 	XG17480 	(g31959,g30673,g4907);
	or 	XG17481 	(g29730,g28141,g28150);
	not 	XG17482 	(g30565,I28832);
	or 	XG17483 	(g33582,g18444,g33351);
	or 	XG17484 	(g32250,g29351,g30598);
	or 	XG17485 	(g30824,g29789,g13833);
	and 	XG17486 	(g32183,g31653,g2795);
	not 	XG17487 	(g29725,g28349);
	not 	XG17488 	(g29697,g28336);
	or 	XG17489 	(g33587,g18463,g33363);
	not 	XG17490 	(I28336,g29147);
	and 	XG17491 	(g32084,g30825,g10948);
	and 	XG17492 	(g32020,g30937,g4157);
	and 	XG17493 	(g31991,g30673,g4912);
	and 	XG17494 	(g32265,g30567,g2799);
	and 	XG17495 	(g32085,g31021,g27253);
	and 	XG17496 	(g32089,g31021,g27261);
	or 	XG17497 	(g32225,g29336,g30576);
	or 	XG17498 	(g33393,g29984,g32286);
	and 	XG17499 	(g32105,g30673,g4922);
	and 	XG17500 	(g32098,g30614,g4732);
	and 	XG17501 	(g32018,g30937,g4146);
	and 	XG17502 	(g31489,g30305,g2204);
	and 	XG17503 	(g32163,g31170,g3502);
	or 	XG17504 	(g29286,g18759,g28542);
	or 	XG17505 	(g30458,g24330,g30005);
	or 	XG17506 	(g32238,g29349,g30594);
	not 	XG17507 	(I29363,g30218);
	and 	XG17508 	(g31273,g27779,g30143);
	and 	XG17509 	(g31296,g27779,g30119);
	and 	XG17510 	(g31282,g27779,g30130);
	and 	XG17511 	(g32170,g27779,g31671);
	and 	XG17512 	(g32042,g31070,g27244);
	and 	XG17513 	(g32055,g30825,g10999);
	and 	XG17514 	(g31513,g29318,g2606);
	or 	XG17515 	(g31871,g18279,g30596);
	or 	XG17516 	(g33588,g18468,g33334);
	and 	XG17517 	(g32287,g30578,g2823);
	or 	XG17518 	(g33598,g18496,g33364);
	and 	XG17519 	(g31501,g29310,g2047);
	and 	XG17520 	(g32278,g30572,g2811);
	or 	XG17521 	(g33276,g29566,g32128);
	or 	XG17522 	(g33590,g18470,g33358);
	or 	XG17523 	(g31869,g18221,g30592);
	or 	XG17524 	(g32230,g29345,g30589);
	and 	XG17525 	(g32070,g30825,g10967);
	or 	XG17526 	(g33579,g18437,g33357);
	and 	XG17527 	(g31323,g27907,g30150);
	or 	XG17528 	(g33270,g29547,g32119);
	and 	XG17529 	(g31283,g27837,g30156);
	and 	XG17530 	(g31297,g27837,g30144);
	or 	XG17531 	(g33580,g18442,g33330);
	or 	XG17532 	(g33589,g18469,g33340);
	or 	XG17533 	(g29257,g18600,g28228);
	not 	XG17534 	(g33426,g32017);
	not 	XG17535 	(I29149,g29384);
	not 	XG17536 	(I27718,g28231);
	or 	XG17537 	(g30984,g29755,g29765);
	not 	XG17538 	(I29139,g29382);
	not 	XG17539 	(I29368,g30321);
	not 	XG17540 	(I27713,g28224);
	and 	XG17541 	(g30269,g23970,g28778);
	and 	XG17542 	(g30284,g23994,g28852);
	and 	XG17543 	(g30235,g23915,g28723);
	and 	XG17544 	(g30216,g23882,g28691);
	and 	XG17545 	(g30194,g23849,g28651);
	and 	XG17546 	(g30226,g23898,g28707);
	and 	XG17547 	(g32010,g22303,g31785);
	and 	XG17548 	(g30257,g23952,g28750);
	and 	XG17549 	(g32009,g22224,g31782);
	and 	XG17550 	(g29347,g22201,g29176);
	and 	XG17551 	(g32305,g20567,g31287);
	and 	XG17552 	(g29326,g22155,g29105);
	and 	XG17553 	(g31967,g22167,g31755);
	and 	XG17554 	(g30166,g23792,g28621);
	and 	XG17555 	(g30230,g23906,g28717);
	and 	XG17556 	(g31986,g22197,g31766);
	and 	XG17557 	(g30198,g23860,g28662);
	and 	XG17558 	(g30178,g23815,g28632);
	and 	XG17559 	(g30188,g23841,g28644);
	and 	XG17560 	(g30154,g23769,g28611);
	and 	XG17561 	(g32273,g20446,g31255);
	and 	XG17562 	(g32301,g20547,g31276);
	and 	XG17563 	(g32306,g23499,g31289);
	and 	XG17564 	(g29806,g23271,g28358);
	and 	XG17565 	(g29805,g23270,g28357);
	and 	XG17566 	(g29842,g23284,g28372);
	and 	XG17567 	(g29857,g23304,g28386);
	and 	XG17568 	(g29872,g23333,g28401);
	and 	XG17569 	(g29749,g23214,g28295);
	and 	XG17570 	(g29766,g23235,g28316);
	and 	XG17571 	(g29871,g23332,g28400);
	and 	XG17572 	(g29757,g23221,g28305);
	and 	XG17573 	(g29783,g23246,g28329);
	and 	XG17574 	(g29747,g23196,g28286);
	and 	XG17575 	(g29794,g23256,g28342);
	and 	XG17576 	(g30001,g23486,g28490);
	and 	XG17577 	(g29758,g23222,g28306);
	and 	XG17578 	(g32324,g23537,g31315);
	and 	XG17579 	(g29841,g23283,g28371);
	and 	XG17580 	(g29856,g23303,g28385);
	and 	XG17581 	(g29885,g23350,g28416);
	and 	XG17582 	(g29782,g23245,g28328);
	and 	XG17583 	(g32323,g20610,g31311);
	and 	XG17584 	(g32291,g20527,g31268);
	and 	XG17585 	(g30191,g23843,g28647);
	and 	XG17586 	(g30211,g23878,g28685);
	and 	XG17587 	(g30190,g23842,g28646);
	and 	XG17588 	(g30199,g23861,g28664);
	and 	XG17589 	(g30223,g23895,g28702);
	and 	XG17590 	(g31968,g22168,g31757);
	and 	XG17591 	(g31976,g22178,g31762);
	and 	XG17592 	(g30210,g23877,g28684);
	and 	XG17593 	(g30233,g23913,g28720);
	and 	XG17594 	(g30272,g23982,g28814);
	and 	XG17595 	(g30200,g23862,g28665);
	and 	XG17596 	(g30180,g23820,g28635);
	and 	XG17597 	(g30243,g23929,g28731);
	and 	XG17598 	(g31987,g22198,g31767);
	and 	XG17599 	(g30254,g23944,g28747);
	and 	XG17600 	(g31237,g25325,g29366);
	and 	XG17601 	(g31242,g25409,g29373);
	and 	XG17602 	(g31996,g18979,g31779);
	and 	XG17603 	(g30219,g23887,g28698);
	and 	XG17604 	(g31966,g22166,g31754);
	and 	XG17605 	(g31974,g22176,g31760);
	and 	XG17606 	(g30248,g23938,g28743);
	and 	XG17607 	(g30208,g23875,g28681);
	and 	XG17608 	(g30140,g23749,g28600);
	and 	XG17609 	(g30207,g23874,g28680);
	and 	XG17610 	(g30175,g23813,g28629);
	and 	XG17611 	(g29320,g22147,g29068);
	and 	XG17612 	(g30165,g23788,g28619);
	and 	XG17613 	(g30228,g23903,g28715);
	and 	XG17614 	(g30152,g23767,g28609);
	and 	XG17615 	(g30196,g23858,g28659);
	and 	XG17616 	(g30239,g23923,g28728);
	and 	XG17617 	(g30186,g23839,g28641);
	and 	XG17618 	(g30185,g23838,g28640);
	and 	XG17619 	(g31960,g22153,g31749);
	and 	XG17620 	(g30238,g23922,g28727);
	and 	XG17621 	(g30229,g23904,g28716);
	and 	XG17622 	(g30164,g23787,g28618);
	and 	XG17623 	(g30153,g23768,g28610);
	and 	XG17624 	(g32269,g20443,g31253);
	and 	XG17625 	(g32330,g20631,g31320);
	and 	XG17626 	(g32300,g20544,g31274);
	and 	XG17627 	(g32256,g20382,g31249);
	and 	XG17628 	(g32241,g20323,g31244);
	and 	XG17629 	(g29899,g23375,g28428);
	and 	XG17630 	(g29875,g23337,g28403);
	and 	XG17631 	(g29874,g23336,g28402);
	and 	XG17632 	(g29843,g23289,g28373);
	and 	XG17633 	(g32332,g23558,g31325);
	and 	XG17634 	(g29770,g23238,g28320);
	and 	XG17635 	(g30024,g23501,g28497);
	and 	XG17636 	(g32307,g23500,g31291);
	and 	XG17637 	(g29784,g23247,g28331);
	and 	XG17638 	(g29807,g23272,g28359);
	and 	XG17639 	(g29759,g23226,g28308);
	and 	XG17640 	(g29795,g23257,g28344);
	and 	XG17641 	(g29859,g23307,g28388);
	and 	XG17642 	(g29751,g23216,g28297);
	and 	XG17643 	(g29887,g23351,g28417);
	and 	XG17644 	(g32314,g23516,g31304);
	and 	XG17645 	(g29785,g23248,g28332);
	and 	XG17646 	(g32322,g20605,g31308);
	and 	XG17647 	(g32242,g20324,g31245);
	and 	XG17648 	(g32292,g20530,g31269);
	and 	XG17649 	(g32312,g20591,g31302);
	and 	XG17650 	(g30267,g23967,g28776);
	and 	XG17651 	(g30266,g23966,g28775);
	and 	XG17652 	(g31993,g22214,g31774);
	and 	XG17653 	(g30275,g23984,g28816);
	and 	XG17654 	(g30203,g23864,g28668);
	and 	XG17655 	(g30234,g23914,g28721);
	and 	XG17656 	(g30245,g23935,g28733);
	and 	XG17657 	(g29337,g22180,g29166);
	and 	XG17658 	(g31977,g22179,g31764);
	and 	XG17659 	(g30246,g23936,g28734);
	and 	XG17660 	(g30281,g23992,g28850);
	and 	XG17661 	(g30274,g23983,g28815);
	and 	XG17662 	(g30192,g23847,g28649);
	and 	XG17663 	(g31988,g22199,g31768);
	and 	XG17664 	(g30225,g23897,g28705);
	and 	XG17665 	(g29797,g23259,g28347);
	and 	XG17666 	(g29798,g23260,g28348);
	and 	XG17667 	(g32333,g23559,g31326);
	and 	XG17668 	(g29861,g23313,g28390);
	and 	XG17669 	(g32326,g23539,g31317);
	and 	XG17670 	(g29808,g23273,g28361);
	and 	XG17671 	(g29845,g23291,g28375);
	and 	XG17672 	(g29909,g23388,g28435);
	and 	XG17673 	(g29788,g23250,g28335);
	and 	XG17674 	(g29876,g23339,g28404);
	and 	XG17675 	(g29772,g23243,g28323);
	and 	XG17676 	(g32315,g23517,g31306);
	and 	XG17677 	(g29809,g23274,g28362);
	and 	XG17678 	(g29787,g23249,g28334);
	and 	XG17679 	(g29891,g23356,g28420);
	and 	XG17680 	(g32304,g20564,g31284);
	and 	XG17681 	(g29987,g22763,g26424,g29197);
	or 	XG17682 	(g33275,g29564,g32127);
	or 	XG17683 	(g33387,g29954,g32263);
	or 	XG17684 	(g33253,g29511,g32103);
	nand 	XG17685 	(g31971,g10511,g30573);
	or 	XG17686 	(g33268,g29538,g32116);
	nand 	XG17687 	(g29540,g13464,g28336);
	or 	XG17688 	(g33257,g29519,g32108);
	nand 	XG17689 	(g31978,g15591,g30580);
	nor 	XG17690 	(g30282,g29073,g6336);
	and 	XG17691 	(g29322,g6336,g7074,g29192);
	nor 	XG17692 	(g30288,g29073,g7087);
	nand 	XG17693 	(g27925,I26440,I26439);
	nor 	XG17694 	(g30276,g29073,g7074);
	and 	XG17695 	(g31300,g27858,g30148);
	and 	XG17696 	(g32175,g27858,g31709);
	and 	XG17697 	(g31286,g27858,g30159);
	and 	XG17698 	(g31312,g27858,g30136);
	and 	XG17699 	(g31275,g27800,g30147);
	and 	XG17700 	(g32171,g27800,g31706);
	and 	XG17701 	(g31299,g27800,g30123);
	and 	XG17702 	(g31285,g27800,g30134);
	nand 	XG17703 	(g31950,g30573,g7285);
	or 	XG17704 	(g33281,g29576,g32142);
	nand 	XG17705 	(g29556,g13486,g28349);
	or 	XG17706 	(g33389,g29964,g32272);
	or 	XG17707 	(g33390,g29968,g32276);
	nor 	XG17708 	(g29903,g28484,g6928);
	and 	XG17709 	(g32178,g27886,g31747);
	and 	XG17710 	(g31321,g27886,g30146);
	and 	XG17711 	(g31310,g27886,g30157);
	and 	XG17712 	(g31298,g27886,g30169);
	and 	XG17713 	(g32174,g27837,g31708);
	and 	XG17714 	(g31309,g27837,g30132);
	nand 	XG17715 	(g31997,g30580,g22306);
	and 	XG17716 	(g31324,g27937,g30171);
	and 	XG17717 	(g31314,g27937,g30183);
	and 	XG17718 	(g32182,g27937,g31753);
	and 	XG17719 	(g31467,g27937,g30162);
	and 	XG17720 	(g31301,g27907,g30170);
	and 	XG17721 	(g32179,g27907,g31748);
	and 	XG17722 	(g31313,g27907,g30160);
	nor 	XG17723 	(g30273,g29036,g5990);
	and 	XG17724 	(g29315,g5990,g7051,g29188);
	nor 	XG17725 	(g30280,g29036,g7064);
	nor 	XG17726 	(g29886,g28458,g3288);
	and 	XG17727 	(g29316,g3288,g6875,g28528);
	nor 	XG17728 	(g29898,g28458,g6895);
	nor 	XG17729 	(g30249,g28982,g5297);
	and 	XG17730 	(g30308,g5297,g7004,g29178);
	nor 	XG17731 	(g30260,g28982,g7018);
	or 	XG17732 	(g33280,g29574,g32141);
	or 	XG17733 	(g33294,g29604,g32152);
	or 	XG17734 	(g33292,g29601,g32150);
	nor 	XG17735 	(g29910,g28484,g3990);
	and 	XG17736 	(g29328,g3990,g6928,g28553);
	nor 	XG17737 	(g29915,g28484,g6941);
	nor 	XG17738 	(g29900,g28471,g3639);
	and 	XG17739 	(g29323,g3639,g6905,g28539);
	nor 	XG17740 	(g29908,g28471,g6918);
	nand 	XG17741 	(g27380,I26072,I26071);
	and 	XG17742 	(g31488,g30302,g1779);
	or 	XG17743 	(g33289,g29588,g32148);
	or 	XG17744 	(g33293,g29602,g32151);
	and 	XG17745 	(g31266,g27742,g30129);
	and 	XG17746 	(g32165,g27742,g31669);
	and 	XG17747 	(g31281,g27742,g30106);
	and 	XG17748 	(g31272,g27742,g30117);
	nand 	XG17749 	(g27955,I26461,I26460);
	not 	XG17750 	(g31667,g30142);
	or 	XG17751 	(g33296,g29617,g32156);
	nand 	XG17752 	(g27767,I26368,I26367);
	nor 	XG17753 	(g30265,g29036,g7051);
	nand 	XG17754 	(g27365,I26051,I26050);
	nor 	XG17755 	(g30240,g28982,g7004);
	or 	XG17756 	(g32427,g30583,g8928);
	nor 	XG17757 	(g30290,g29110,g6682);
	and 	XG17758 	(g30316,g6682,g7097,g29199);
	nor 	XG17759 	(g30294,g29110,g7110);
	nand 	XG17760 	(g27824,I26395,I26394);
	or 	XG17761 	(g33262,g29528,g32112);
	nor 	XG17762 	(g30285,g29110,g7097);
	or 	XG17763 	(g33261,g29525,g32111);
	nand 	XG17764 	(g27876,I26419,I26418);
	nand 	XG17765 	(g27401,I26095,I26094);
	nor 	XG17766 	(g29889,g28471,g6905);
	or 	XG17767 	(g33260,g29524,g32110);
	or 	XG17768 	(g32408,g30073,g31541);
	or 	XG17769 	(g33571,g18409,g33367);
	nor 	XG17770 	(g31970,g30583,g9024);
	nor 	XG17771 	(g31965,g4358,g30583);
	or 	XG17772 	(g33604,g18520,g33345);
	or 	XG17773 	(g33550,g18338,g33342);
	or 	XG17774 	(g33556,g18362,g33329);
	nor 	XG17775 	(g31942,g30583,g8977);
	nor 	XG17776 	(g31935,g4349,g30583);
	or 	XG17777 	(g29263,g18617,g28239);
	or 	XG17778 	(g33573,g18415,g33343);
	or 	XG17779 	(g33606,g18522,g33369);
	or 	XG17780 	(g29280,g18742,g28530);
	or 	XG17781 	(g33565,g18389,g33338);
	or 	XG17782 	(g33572,g18414,g33339);
	or 	XG17783 	(g33603,g18515,g33372);
	or 	XG17784 	(g33558,g18364,g33350);
	not 	XG17785 	(g34351,g34174);
	or 	XG17786 	(g33605,g18521,g33352);
	nand 	XG17787 	(g33669,g862,g33378);
	or 	XG17788 	(g33557,g18363,g33331);
	or 	XG17789 	(g33548,g18336,g33327);
	or 	XG17790 	(g33555,g18357,g33355);
	or 	XG17791 	(g33960,g21701,g33759);
	not 	XG17792 	(g33250,g32186);
	or 	XG17793 	(g33574,g18416,g33362);
	or 	XG17794 	(g33547,g18331,g33349);
	or 	XG17795 	(g33549,g18337,g33328);
	or 	XG17796 	(g32398,g30061,g31526);
	or 	XG17797 	(g29269,g18634,g28249);
	or 	XG17798 	(g33564,g18388,g33332);
	or 	XG17799 	(g29292,g18776,g28556);
	and 	XG17800 	(g30278,g23988,g28818);
	and 	XG17801 	(g30205,g23869,g28671);
	and 	XG17802 	(g30204,g23868,g28670);
	and 	XG17803 	(g30289,g24000,g28884);
	and 	XG17804 	(g30227,g23899,g28708);
	and 	XG17805 	(g30277,g23987,g28817);
	and 	XG17806 	(g30268,g23969,g28777);
	and 	XG17807 	(g30236,g23916,g28724);
	and 	XG17808 	(g30283,g23993,g28851);
	and 	XG17809 	(g30247,g23937,g28735);
	and 	XG17810 	(g30258,g23953,g28751);
	and 	XG17811 	(g30215,g23881,g28690);
	and 	XG17812 	(g32338,g20668,g31466);
	and 	XG17813 	(g32283,g20506,g31259);
	and 	XG17814 	(g32274,g20447,g31256);
	and 	XG17815 	(g30221,g23893,g28700);
	and 	XG17816 	(g30250,g23939,g28744);
	and 	XG17817 	(g30231,g23907,g28718);
	and 	XG17818 	(g30251,g23940,g28745);
	and 	XG17819 	(g30242,g23927,g28730);
	and 	XG17820 	(g30241,g23926,g28729);
	and 	XG17821 	(g30197,g23859,g28661);
	and 	XG17822 	(g30222,g23894,g28701);
	and 	XG17823 	(g30209,g23876,g28682);
	and 	XG17824 	(g30177,g23814,g28631);
	and 	XG17825 	(g30187,g23840,g28643);
	and 	XG17826 	(g30261,g23961,g28772);
	and 	XG17827 	(g30167,g23793,g28622);
	and 	XG17828 	(g32261,g20386,g31251);
	and 	XG17829 	(g32331,g20637,g31322);
	and 	XG17830 	(g29750,g23215,g28296);
	and 	XG17831 	(g29767,g23236,g28317);
	and 	XG17832 	(g32246,g20326,g31246);
	and 	XG17833 	(g32260,g20385,g31250);
	and 	XG17834 	(g30264,g23963,g28774);
	and 	XG17835 	(g30263,g23962,g28773);
	and 	XG17836 	(g30168,g23794,g28623);
	and 	XG17837 	(g29331,g22169,g29143);
	and 	XG17838 	(g30253,g23943,g28746);
	and 	XG17839 	(g30179,g23819,g28634);
	and 	XG17840 	(g30244,g23930,g28732);
	and 	XG17841 	(g30232,g23912,g28719);
	and 	XG17842 	(g30174,g23812,g28628);
	and 	XG17843 	(g30220,g23888,g28699);
	and 	XG17844 	(g31990,g18945,g31772);
	and 	XG17845 	(g29796,g23258,g28345);
	and 	XG17846 	(g29888,g23352,g28418);
	and 	XG17847 	(g29760,g23227,g28309);
	and 	XG17848 	(g29844,g23290,g28374);
	and 	XG17849 	(g29858,g23306,g28387);
	and 	XG17850 	(g29769,g23237,g28319);
	and 	XG17851 	(g32343,g20710,g31473);
	and 	XG17852 	(g32284,g20507,g31260);
	and 	XG17853 	(g34348,g20128,g34125);
	and 	XG17854 	(g34146,g20091,g33788);
	and 	XG17855 	(g30212,g23879,g28687);
	and 	XG17856 	(g30193,g23848,g28650);
	and 	XG17857 	(g30256,g23947,g28749);
	and 	XG17858 	(g30255,g23946,g28748);
	and 	XG17859 	(g30202,g23863,g28667);
	and 	XG17860 	(g30181,g23821,g28636);
	and 	XG17861 	(g30224,g23896,g28704);
	and 	XG17862 	(g30213,g23880,g28688);
	and 	XG17863 	(g30041,g23518,g28511);
	and 	XG17864 	(g29860,g23312,g28389);
	and 	XG17865 	(g29890,g23355,g28419);
	and 	XG17866 	(g29902,g23377,g28430);
	and 	XG17867 	(g29901,g23376,g28429);
	and 	XG17868 	(g29771,g23242,g28322);
	and 	XG17869 	(g29877,g23340,g28405);
	and 	XG17870 	(g29761,g23228,g28310);
	and 	XG17871 	(g34322,g34174,g14188);
	nor 	XG17872 	(g34359,g12259,g34174,g9162);
	and 	XG17873 	(g34324,g34161,g14064);
	or 	XG17874 	(g34332,g33723,g34071);
	or 	XG17875 	(g33566,g18390,g33356);
	or 	XG17876 	(g29304,g18810,g28588);
	or 	XG17877 	(g34022,g18538,g33873);
	and 	XG17878 	(g34069,g33797,g8774);
	or 	XG17879 	(g34251,g18147,g34157);
	or 	XG17880 	(g33563,g18383,g33361);
	or 	XG17881 	(g29298,g18793,g28571);
	or 	XG17882 	(g29222,g18105,g28252);
	or 	XG17883 	(g33965,g18179,g33805);
	and 	XG17884 	(g34110,g22935,g33732);
	and 	XG17885 	(g34111,g22936,g33733);
	or 	XG17886 	(g33961,g21712,g33789);
	or 	XG17887 	(g34107,g33121,g33710);
	not 	XG17888 	(g34147,g33823);
	and 	XG17889 	(g34073,g33823,g8948);
	nand 	XG17890 	(g34162,g11679,g33823,g785);
	and 	XG17891 	(g32187,g25287,g30672);
	and 	XG17892 	(g32194,g28436,g30601);
	not 	XG17893 	(I29199,g30237);
	not 	XG17894 	(g32394,g30601);
	not 	XG17895 	(g29041,I27385);
	not 	XG17896 	(I29977,g31596);
	not 	XG17897 	(g32446,g31596);
	not 	XG17898 	(g32318,g31596);
	nor 	XG17899 	(g33134,g32057,g7686);
	nor 	XG17900 	(g33131,g32057,g4659);
	and 	XG17901 	(g32205,g28463,g30922);
	or 	XG17902 	(g32990,g18341,g32281);
	not 	XG17903 	(g28155,I26664);
	nand 	XG17904 	(g33083,g32118,g7805);
	or 	XG17905 	(I30761,g32082,g32067,g32167,g32071);
	not 	XG17906 	(g30182,I28419);
	or 	XG17907 	(g33001,g18404,g32282);
	not 	XG17908 	(g28142,I26649);
	or 	XG17909 	(g33000,g18403,g32270);
	or 	XG17910 	(g32988,g18325,g32232);
	not 	XG17911 	(g28166,I26687);
	not 	XG17912 	(g28162,I26679);
	or 	XG17913 	(g32994,g18367,g32290);
	not 	XG17914 	(g29491,I27777);
	not 	XG17915 	(g28157,I26670);
	or 	XG17916 	(I30734,g32095,g32086,g32191,g31790);
	not 	XG17917 	(I28349,g28367);
	nor 	XG17918 	(g33141,g8400,g32099);
	not 	XG17919 	(g28262,I26785);
	and 	XG17920 	(g33441,g29722,g32251);
	not 	XG17921 	(g29498,I27784);
	not 	XG17922 	(I27749,g28917);
	or 	XG17923 	(g32999,g18401,g32337);
	and 	XG17924 	(g33429,g29676,g32231);
	and 	XG17925 	(g33450,g29737,g32266);
	not 	XG17926 	(I29582,g30591);
	or 	XG17927 	(I30750,g32070,g32054,g32310,g31788);
	not 	XG17928 	(g28819,I27271);
	or 	XG17929 	(I30718,g32020,g32097,g32356,g32348);
	or 	XG17930 	(I30746,g32309,g31991,g31985,g32047);
	or 	XG17931 	(I30741,g32013,g32224,g32030,g32085);
	or 	XG17932 	(I30735,g32035,g32089,g32376,g32369);
	not 	XG17933 	(g30328,I28585);
	and 	XG17934 	(g31261,g30259,g14754);
	and 	XG17935 	(g31240,g30206,g14793);
	or 	XG17936 	(I30728,g32018,g32056,g32350,g32345);
	or 	XG17937 	(I30756,g32105,g32098,g32163,g32088);
	not 	XG17938 	(g28161,I26676);
	not 	XG17939 	(g33136,g32057);
	not 	XG17940 	(I29913,g30605);
	or 	XG17941 	(I30751,g31959,g31943,g32161,g32042);
	or 	XG17942 	(g33068,g22112,g31994);
	not 	XG17943 	(I27735,g28779);
	and 	XG17944 	(I31122,g32634,g32633,g32632,g32631);
	and 	XG17945 	(I31142,g32664,g32663,g32662,g32661);
	and 	XG17946 	(I31117,g32627,g32626,g32625,g32624);
	and 	XG17947 	(I31087,g32583,g32582,g32581,g32580);
	and 	XG17948 	(I31017,g32483,g32482,g32481,g32480);
	and 	XG17949 	(I31097,g32599,g32598,g32597,g32596);
	and 	XG17950 	(I31032,g32504,g32503,g32502,g32501);
	and 	XG17951 	(I31052,g32534,g32533,g32532,g32531);
	and 	XG17952 	(I31137,g32657,g32656,g32655,g32654);
	and 	XG17953 	(I31127,g32641,g32640,g32639,g32638);
	and 	XG17954 	(I31042,g32518,g32517,g32516,g32515);
	and 	XG17955 	(I31177,g32713,g32712,g32711,g32710);
	and 	XG17956 	(I31037,g32511,g32510,g32509,g32508);
	and 	XG17957 	(I31082,g32576,g32575,g32574,g32573);
	and 	XG17958 	(I31132,g32648,g32647,g32646,g32645);
	and 	XG17959 	(I31102,g32606,g32605,g32604,g32603);
	and 	XG17960 	(I31162,g32692,g32691,g32690,g32689);
	and 	XG17961 	(I31167,g32699,g32698,g32697,g32696);
	and 	XG17962 	(I31002,g32462,g32461,g32460,g32459);
	and 	XG17963 	(I31062,g32548,g32547,g32546,g32545);
	and 	XG17964 	(I31027,g32497,g32496,g32495,g32494);
	and 	XG17965 	(I31147,g32671,g32670,g32669,g32668);
	and 	XG17966 	(I31107,g32613,g32612,g32611,g32610);
	and 	XG17967 	(I31092,g32592,g32591,g32590,g32589);
	and 	XG17968 	(I31047,g32527,g32526,g32525,g32524);
	and 	XG17969 	(I31172,g32706,g32705,g32704,g32703);
	and 	XG17970 	(I31007,g32469,g32468,g32467,g32466);
	and 	XG17971 	(I31072,g32562,g32561,g32560,g32559);
	and 	XG17972 	(I31077,g32569,g32568,g32567,g32566);
	and 	XG17973 	(I31152,g32678,g32677,g32676,g32675);
	and 	XG17974 	(I31057,g32541,g32540,g32539,g32538);
	and 	XG17975 	(I31012,g32476,g32475,g32474,g32473);
	and 	XG17976 	(I31327,g32931,g32930,g32929,g32928);
	and 	XG17977 	(I31237,g32801,g32800,g32799,g32798);
	and 	XG17978 	(I31317,g32917,g32916,g32915,g32914);
	and 	XG17979 	(I31247,g32815,g32814,g32813,g32812);
	and 	XG17980 	(I31342,g32952,g32951,g32950,g32949);
	and 	XG17981 	(I31202,g32750,g32749,g32748,g32747);
	and 	XG17982 	(I31207,g32757,g32756,g32755,g32754);
	and 	XG17983 	(I31227,g32787,g32786,g32785,g32784);
	and 	XG17984 	(I31197,g32743,g32742,g32741,g32740);
	and 	XG17985 	(I31337,g32945,g32944,g32943,g32942);
	and 	XG17986 	(I31272,g32852,g32851,g32850,g32849);
	and 	XG17987 	(I31347,g32959,g32958,g32957,g32956);
	and 	XG17988 	(I31277,g32859,g32858,g32857,g32856);
	and 	XG17989 	(I31182,g32722,g32721,g32720,g32719);
	and 	XG17990 	(I31322,g32924,g32923,g32922,g32921);
	and 	XG17991 	(I31192,g32736,g32735,g32734,g32733);
	and 	XG17992 	(I31212,g32764,g32763,g32762,g32761);
	and 	XG17993 	(I31292,g32880,g32879,g32878,g32877);
	and 	XG17994 	(I31302,g32894,g32893,g32892,g32891);
	and 	XG17995 	(I31332,g32938,g32937,g32936,g32935);
	and 	XG17996 	(I31252,g32822,g32821,g32820,g32819);
	and 	XG17997 	(I31282,g32866,g32865,g32864,g32863);
	and 	XG17998 	(I31307,g32901,g32900,g32899,g32898);
	and 	XG17999 	(I31242,g32808,g32807,g32806,g32805);
	and 	XG18000 	(I31312,g32908,g32907,g32906,g32905);
	and 	XG18001 	(I31187,g32729,g32728,g32727,g32726);
	and 	XG18002 	(I31257,g32829,g32828,g32827,g32826);
	and 	XG18003 	(I31232,g32794,g32793,g32792,g32791);
	and 	XG18004 	(I31287,g32873,g32872,g32871,g32870);
	and 	XG18005 	(I31297,g32887,g32886,g32885,g32884);
	and 	XG18006 	(I31222,g32778,g32777,g32776,g32775);
	and 	XG18007 	(I31267,g32843,g32842,g32841,g32840);
	and 	XG18008 	(I31352,g32966,g32965,g32964,g32963);
	and 	XG18009 	(I31262,g32836,g32835,g32834,g32833);
	and 	XG18010 	(I31357,g32973,g32972,g32971,g32970);
	and 	XG18011 	(I31217,g32771,g32770,g32769,g32768);
	nor 	XG18012 	(g32520,I30055,I30054,g31554);
	nor 	XG18013 	(g32455,I29986,I29985,g31566);
	and 	XG18014 	(I31157,g32685,g32684,g32683,g32682);
	nor 	XG18015 	(g32585,I30124,I30123,g31542);
	nor 	XG18016 	(g32650,I30193,I30192,g31579);
	and 	XG18017 	(I31067,g32555,g32554,g32553,g32552);
	and 	XG18018 	(I31022,g32490,g32489,g32488,g32487);
	and 	XG18019 	(I31112,g32620,g32619,g32618,g32617);
	nor 	XG18020 	(g32715,I30262,I30261,g31327);
	nor 	XG18021 	(g32910,I30469,I30468,g31327);
	nor 	XG18022 	(g32780,I30331,I30330,g31327);
	not 	XG18023 	(I27730,g28752);
	not 	XG18024 	(g28184,I26705);
	or 	XG18025 	(I30755,g32055,g32049,g32303,g30564);
	not 	XG18026 	(I28838,g29372);
	or 	XG18027 	(g33034,g21844,g32340);
	not 	XG18028 	(I28301,g29042);
	or 	XG18029 	(I30727,g31941,g31933,g32196,g31759);
	or 	XG18030 	(g33067,g22111,g31989);
	or 	XG18031 	(g33047,g21927,g31944);
	or 	XG18032 	(g33060,g22022,g31992);
	not 	XG18033 	(g28163,I26682);
	nor 	XG18034 	(g32845,I30400,I30399,g30673);
	not 	XG18035 	(I29894,g31771);
	or 	XG18036 	(g33054,g21975,g31975);
	or 	XG18037 	(g31895,g24296,g31505);
	or 	XG18038 	(g33028,g21797,g32325);
	or 	XG18039 	(g33052,g21973,g31961);
	or 	XG18040 	(g32987,g18323,g32311);
	or 	XG18041 	(g32993,g18352,g32255);
	or 	XG18042 	(I30745,g32084,g32069,g32321,g31777);
	not 	XG18043 	(g29185,I27481);
	not 	XG18044 	(g28173,I26693);
	not 	XG18045 	(g28181,I26700);
	not 	XG18046 	(I28540,g28954);
	or 	XG18047 	(g33023,g21751,g32313);
	or 	XG18048 	(g33021,g21749,g32302);
	or 	XG18049 	(g33065,g22068,g32008);
	not 	XG18050 	(g33385,g32038);
	not 	XG18051 	(g33382,g32033);
	and 	XG18052 	(g33886,g20614,g33297);
	and 	XG18053 	(g33863,g20505,g33273);
	and 	XG18054 	(g33872,g20548,g33282);
	and 	XG18055 	(g33884,g20590,g33295);
	and 	XG18056 	(g33857,g20445,g33267);
	and 	XG18057 	(g33866,g20528,g33276);
	and 	XG18058 	(g33841,g20268,g33254);
	and 	XG18059 	(g33878,g20565,g33288);
	and 	XG18060 	(g33943,g21609,g33384);
	and 	XG18061 	(g33862,g20504,g33272);
	and 	XG18062 	(g32184,g25249,g30611);
	and 	XG18063 	(g32189,g25369,g30824);
	and 	XG18064 	(g32164,g25171,g30733);
	and 	XG18065 	(g32206,g25524,g30609);
	and 	XG18066 	(g32168,g25185,g30597);
	and 	XG18067 	(g32177,g25214,g30608);
	and 	XG18068 	(g32199,g25506,g30916);
	and 	XG18069 	(g32195,g25451,g30734);
	and 	XG18070 	(g32193,g25410,g30732);
	and 	XG18071 	(g33856,g20442,g33266);
	and 	XG18072 	(g33639,g18829,g33386);
	and 	XG18073 	(g33843,g20325,g33256);
	and 	XG18074 	(g33877,g20563,g33287);
	and 	XG18075 	(g33941,g21560,g33380);
	and 	XG18076 	(g33868,g20542,g33278);
	and 	XG18077 	(g33837,g20233,g33251);
	and 	XG18078 	(g33842,g20322,g33255);
	and 	XG18079 	(g33864,g20524,g33274);
	and 	XG18080 	(g33855,g20441,g33265);
	and 	XG18081 	(g33869,g20543,g33279);
	and 	XG18082 	(g33942,g21608,g33383);
	and 	XG18083 	(g33846,g20380,g33259);
	and 	XG18084 	(g33860,g20501,g33270);
	and 	XG18085 	(g33876,g20562,g33286);
	and 	XG18086 	(g33880,g20568,g33290);
	and 	XG18087 	(g33887,g20615,g33298);
	and 	XG18088 	(g33889,g20641,g33303);
	and 	XG18089 	(g33867,g20529,g33277);
	and 	XG18090 	(g33652,g18889,g33393);
	and 	XG18091 	(g33861,g20502,g33271);
	not 	XG18092 	(g29353,I27713);
	not 	XG18093 	(g31794,I29368);
	not 	XG18094 	(g31479,I29139);
	not 	XG18095 	(I29961,g30984);
	not 	XG18096 	(g32430,g30984);
	not 	XG18097 	(g32377,g30984);
	not 	XG18098 	(g29358,I27718);
	not 	XG18099 	(g31487,I29149);
	and 	XG18100 	(I31271,g32848,g32847,g32846,g29385);
	and 	XG18101 	(I31316,g32913,g32912,g32911,g29385);
	and 	XG18102 	(I31046,g32523,g32522,g32521,g29385);
	and 	XG18103 	(I31091,g32588,g32587,g32586,g29385);
	and 	XG18104 	(I31136,g32653,g32652,g32651,g29385);
	and 	XG18105 	(I31001,g32458,g32457,g32456,g29385);
	and 	XG18106 	(I31181,g32718,g32717,g32716,g29385);
	and 	XG18107 	(I31226,g32783,g32782,g32781,g29385);
	and 	XG18108 	(I31296,g32883,g32882,g31848,g30937);
	and 	XG18109 	(I31301,g32890,g32889,g31849,g31327);
	and 	XG18110 	(I31056,g32537,g32536,g31805,g30735);
	and 	XG18111 	(I31016,g32479,g32478,g31798,g30825);
	and 	XG18112 	(I31101,g32602,g32601,g31813,g30735);
	and 	XG18113 	(I31021,g32486,g32485,g31799,g31070);
	and 	XG18114 	(I31321,g32920,g32919,g31852,g31376);
	and 	XG18115 	(I31071,g32558,g32557,g31808,g31170);
	and 	XG18116 	(I31076,g32565,g32564,g31809,g30614);
	and 	XG18117 	(I31231,g32790,g32789,g31836,g31376);
	and 	XG18118 	(I31326,g32927,g32926,g31853,g30735);
	and 	XG18119 	(I31151,g32674,g32673,g31822,g30825);
	and 	XG18120 	(I31236,g32797,g32796,g31837,g30735);
	and 	XG18121 	(I31196,g32739,g32738,g31830,g30825);
	and 	XG18122 	(I31261,g32832,g32831,g31842,g30937);
	and 	XG18123 	(I31116,g32623,g32622,g31816,g31154);
	and 	XG18124 	(I31156,g32681,g32680,g31823,g31070);
	and 	XG18125 	(I31121,g32630,g32629,g31817,g30614);
	and 	XG18126 	(I31081,g32572,g32571,g31810,g30673);
	and 	XG18127 	(I31266,g32839,g32838,g31843,g31327);
	and 	XG18128 	(I31201,g32746,g32745,g31831,g31672);
	and 	XG18129 	(I31341,g32948,g32947,g31856,g31710);
	and 	XG18130 	(I31346,g32955,g32954,g31857,g31021);
	and 	XG18131 	(I31036,g32507,g32506,g31802,g30673);
	and 	XG18132 	(I31306,g32897,g32896,g31850,g30614);
	and 	XG18133 	(I31086,g32579,g32578,g31811,g31554);
	and 	XG18134 	(I31171,g32702,g32701,g31826,g31528);
	and 	XG18135 	(I31041,g32514,g32513,g31803,g31566);
	and 	XG18136 	(I31176,g32709,g32708,g31827,g31579);
	and 	XG18137 	(I31286,g32869,g32868,g31846,g30825);
	and 	XG18138 	(I31141,g32660,g32659,g31820,g31376);
	and 	XG18139 	(I31311,g32904,g32903,g31851,g30673);
	and 	XG18140 	(I31291,g32876,g32875,g31847,g31021);
	and 	XG18141 	(I31251,g32818,g32817,g31840,g31710);
	and 	XG18142 	(I31006,g32465,g32464,g31796,g31376);
	and 	XG18143 	(I31011,g32472,g32471,g31797,g30735);
	and 	XG18144 	(I31216,g32767,g32766,g31834,g30937);
	and 	XG18145 	(I31146,g32667,g32666,g31821,g30735);
	and 	XG18146 	(I31061,g32544,g32543,g31806,g30825);
	and 	XG18147 	(I31221,g32774,g32773,g31835,g31327);
	and 	XG18148 	(I31256,g32825,g32824,g31841,g31021);
	and 	XG18149 	(I31066,g32551,g32550,g31807,g31070);
	and 	XG18150 	(I31106,g32609,g32608,g31814,g30825);
	and 	XG18151 	(I31026,g32493,g32492,g31800,g31194);
	and 	XG18152 	(I31111,g32616,g32615,g31815,g31070);
	and 	XG18153 	(I31241,g32804,g32803,g31838,g30825);
	and 	XG18154 	(I31246,g32811,g32810,g31839,g31672);
	and 	XG18155 	(I31331,g32934,g32933,g31854,g30825);
	and 	XG18156 	(I31031,g32500,g32499,g31801,g30614);
	and 	XG18157 	(I31126,g32637,g32636,g31818,g30673);
	and 	XG18158 	(I31131,g32644,g32643,g31819,g31542);
	and 	XG18159 	(I31336,g32941,g32940,g31855,g31672);
	and 	XG18160 	(I31161,g32688,g32687,g31824,g30614);
	and 	XG18161 	(I31276,g32855,g32854,g31844,g31376);
	and 	XG18162 	(I31351,g32962,g32961,g31858,g30937);
	and 	XG18163 	(I31166,g32695,g32694,g31825,g30673);
	and 	XG18164 	(I31356,g32969,g32968,g31859,g31327);
	and 	XG18165 	(I31206,g32753,g32752,g31832,g31710);
	and 	XG18166 	(I31281,g32862,g32861,g31845,g30735);
	and 	XG18167 	(I31186,g32725,g32724,g31828,g31376);
	and 	XG18168 	(I31191,g32732,g32731,g31829,g30735);
	and 	XG18169 	(I31096,g32595,g32594,g31812,g31376);
	and 	XG18170 	(I31211,g32760,g32759,g31833,g31021);
	and 	XG18171 	(I31051,g32530,g32529,g31804,g31376);
	or 	XG18172 	(g32426,g30613,g26131,g26105);
	or 	XG18173 	(g32357,g31296,g29865);
	and 	XG18174 	(g31207,g20739,g30252);
	nor 	XG18175 	(g33147,g7788,g32090);
	or 	XG18176 	(g32353,g31283,g29853);
	and 	XG18177 	(g30914,g20887,g29873);
	nor 	XG18178 	(g33163,g7809,g32099);
	nor 	XG18179 	(g33175,g7828,g32099);
	or 	XG18180 	(I30717,g31949,g31940,g32200,g31787);
	nor 	XG18181 	(g33128,g32057,g4653);
	nor 	XG18182 	(g33125,g32057,g8606);
	or 	XG18183 	(g32347,g31273,g29839);
	and 	XG18184 	(g31936,g24005,g31213);
	and 	XG18185 	(g33440,g29719,g32250);
	and 	XG18186 	(g33423,g29657,g32225);
	or 	XG18187 	(g33312,g32170,g29646);
	or 	XG18188 	(I29352,g30308,g30315,g29315,g29322);
	nor 	XG18189 	(g33144,g32057,g4664);
	nor 	XG18190 	(g33139,g32057,g8650);
	nor 	XG18191 	(g33133,g31503,g32278);
	or 	XG18192 	(g32390,g29979,g31501);
	or 	XG18193 	(g29914,I28147,g22585,g22531);
	or 	XG18194 	(g32352,g31282,g29852);
	or 	XG18195 	(g32392,g30000,g31513);
	or 	XG18196 	(I30760,g32050,g32046,g32295,g31778);
	nor 	XG18197 	(g33138,g31514,g32287);
	nor 	XG18198 	(g33146,g32057,g4669);
	nor 	XG18199 	(g33160,g32057,g8672);
	and 	XG18200 	(g31969,g22139,g31189);
	or 	XG18201 	(g32388,g29962,g31495);
	not 	XG18202 	(g31791,I29363);
	or 	XG18203 	(g32385,g29938,g31480);
	or 	XG18204 	(g32387,g29952,g31489);
	nor 	XG18205 	(g33161,g7806,g32090);
	nor 	XG18206 	(g33130,g31497,g32265);
	nor 	XG18207 	(g33135,g8350,g32090);
	not 	XG18208 	(g30105,I28336);
	nor 	XG18209 	(g33108,g31228,g32183);
	not 	XG18210 	(I29579,g30565);
	not 	XG18211 	(I28866,g29730);
	or 	XG18212 	(g32391,g29982,g31502);
	and 	XG18213 	(g33434,g29702,g32239);
	and 	XG18214 	(g32336,g11842,g31596);
	or 	XG18215 	(g32389,g29966,g31496);
	nor 	XG18216 	(g33107,g31223,g32180);
	nor 	XG18217 	(g33148,g32072,g4854);
	nor 	XG18218 	(g33145,g32072,g8677);
	nor 	XG18219 	(g33137,g32072,g4849);
	not 	XG18220 	(g33142,g32072);
	nor 	XG18221 	(g33100,g31188,g32172);
	not 	XG18222 	(g32421,g31213);
	not 	XG18223 	(I29973,g31213);
	not 	XG18224 	(g32442,g31213);
	nor 	XG18225 	(g33143,g31518,g32293);
	nor 	XG18226 	(g33103,g31212,g32176);
	not 	XG18227 	(g32434,g31189);
	not 	XG18228 	(g31945,g31189);
	not 	XG18229 	(I29965,g31189);
	not 	XG18230 	(g32329,g31522);
	and 	XG18231 	(g31218,g23909,g30271);
	and 	XG18232 	(g31208,g25188,g30262);
	or 	XG18233 	(I30740,g32087,g32083,g32188,g31776);
	not 	XG18234 	(g32393,g30922);
	or 	XG18235 	(g32359,g31298,g29867);
	nor 	XG18236 	(g33427,g31950,g10278);
	nor 	XG18237 	(g33097,g4628,g31950);
	or 	XG18238 	(g30411,g21770,g29872);
	or 	XG18239 	(g33029,g21798,g32332);
	or 	XG18240 	(g30477,g21948,g30239);
	or 	XG18241 	(g30404,g21763,g29758);
	or 	XG18242 	(g30399,g21758,g29757);
	nor 	XG18243 	(g33419,g7627,g31978);
	nor 	XG18244 	(g33085,g4311,g31978);
	or 	XG18245 	(g30398,g21757,g29749);
	or 	XG18246 	(g33316,g32178,g29685);
	or 	XG18247 	(g30539,g22085,g30267);
	or 	XG18248 	(g30397,g21756,g29747);
	or 	XG18249 	(g30441,g21850,g29787);
	and 	XG18250 	(g30915,g24778,g29886);
	and 	XG18251 	(g30919,g23286,g29898);
	or 	XG18252 	(g33009,g18458,g32273);
	nor 	XG18253 	(g33129,g32072,g8630);
	nor 	XG18254 	(g33132,g32072,g4843);
	or 	XG18255 	(g30465,g21936,g30164);
	and 	XG18256 	(g30921,g24789,g29900);
	and 	XG18257 	(g30925,g23309,g29908);
	or 	XG18258 	(g30540,g22086,g30275);
	or 	XG18259 	(g33048,g21928,g31960);
	or 	XG18260 	(g30554,g22125,g30216);
	or 	XG18261 	(g30507,g22028,g30190);
	or 	XG18262 	(g30412,g21771,g29885);
	or 	XG18263 	(g33069,g22113,g32009);
	or 	XG18264 	(g30395,g21754,g29841);
	or 	XG18265 	(g30421,g21805,g29784);
	or 	XG18266 	(g30430,g21814,g29859);
	or 	XG18267 	(g33002,g18419,g32304);
	or 	XG18268 	(g32370,g31312,g29882);
	or 	XG18269 	(g32986,g18280,g31996);
	or 	XG18270 	(g30402,g21761,g29871);
	or 	XG18271 	(g30474,g21945,g30208);
	or 	XG18272 	(g30413,g21772,g30001);
	or 	XG18273 	(g30401,g21760,g29782);
	or 	XG18274 	(g32995,g18375,g32330);
	nor 	XG18275 	(g31469,g29725,g8822);
	nor 	XG18276 	(g31373,g29725,g4975);
	or 	XG18277 	(g30400,g21759,g29766);
	or 	XG18278 	(g30469,g21940,g30153);
	or 	XG18279 	(g30434,g21818,g30024);
	or 	XG18280 	(g30551,g22122,g30235);
	or 	XG18281 	(g30450,g21859,g29861);
	or 	XG18282 	(g33070,g22114,g32010);
	or 	XG18283 	(g32362,g31301,g29870);
	or 	XG18284 	(g32354,g31285,g29854);
	or 	XG18285 	(g30445,g21854,g29772);
	or 	XG18286 	(g32346,g31272,g29838);
	or 	XG18287 	(g30541,g22087,g30281);
	or 	XG18288 	(g33317,g32179,g29688);
	nor 	XG18289 	(g33174,g32072,g8714);
	nor 	XG18290 	(g33162,g32072,g4859);
	or 	XG18291 	(g33049,g21929,g31966);
	or 	XG18292 	(g30516,g22037,g30233);
	nor 	XG18293 	(g33447,g7643,g31978);
	nor 	XG18294 	(g33089,g4322,g31978);
	or 	XG18295 	(g30544,g22115,g30257);
	or 	XG18296 	(g32997,g18378,g32269);
	or 	XG18297 	(g30511,g22032,g30180);
	or 	XG18298 	(g32344,g31266,g29804);
	or 	XG18299 	(g32360,g31299,g29868);
	or 	XG18300 	(g30462,g21933,g30228);
	nor 	XG18301 	(g33140,g32072,g7693);
	or 	XG18302 	(g30547,g22118,g30194);
	or 	XG18303 	(g30531,g22077,g30274);
	or 	XG18304 	(g32361,g31300,g29869);
	or 	XG18305 	(g32373,g31321,g29894);
	or 	XG18306 	(g30446,g21855,g29788);
	or 	XG18307 	(g32991,g18349,g32322);
	or 	XG18308 	(g30471,g21942,g30175);
	or 	XG18309 	(g33053,g21974,g31967);
	and 	XG18310 	(g31231,g25239,g30290);
	and 	XG18311 	(g31232,g23972,g30294);
	or 	XG18312 	(g30473,g21944,g30196);
	or 	XG18313 	(g30452,g21861,g29891);
	or 	XG18314 	(g33062,g22065,g31977);
	or 	XG18315 	(g30468,g21939,g30238);
	or 	XG18316 	(g30512,g22033,g30191);
	or 	XG18317 	(g30447,g21856,g29798);
	or 	XG18318 	(g30523,g22069,g30245);
	nor 	XG18319 	(g31133,g29556,g7953);
	nor 	XG18320 	(g31127,g29556,g4966);
	or 	XG18321 	(g33055,g21976,g31986);
	or 	XG18322 	(g30536,g22082,g30234);
	or 	XG18323 	(g30492,g21988,g30188);
	nor 	XG18324 	(g31372,g29697,g8796);
	nor 	XG18325 	(g31318,g29697,g4785);
	nor 	XG18326 	(g31491,g29725,g8938);
	nor 	XG18327 	(g31483,g29725,g4899);
	or 	XG18328 	(g33006,g18447,g32291);
	or 	XG18329 	(g32374,g31323,g29895);
	or 	XG18330 	(I29351,g30316,g29316,g29323,g29328);
	or 	XG18331 	(g30518,g22039,g30254);
	or 	XG18332 	(g30449,g21858,g29845);
	or 	XG18333 	(g30513,g22034,g30200);
	and 	XG18334 	(g33304,g31971,g32427);
	and 	XG18335 	(g33859,g10531,g33426);
	nor 	XG18336 	(g31482,g29697,g8883);
	and 	XG18337 	(g33428,g29672,g32230);
	nor 	XG18338 	(g31476,g29697,g4709);
	and 	XG18339 	(g33433,g29694,g32238);
	nor 	XG18340 	(g31119,g29556,g7898);
	nor 	XG18341 	(g31117,g29556,g4991);
	and 	XG18342 	(g31183,g25174,g30249);
	and 	XG18343 	(g31206,g23890,g30260);
	and 	XG18344 	(g31220,g25202,g30273);
	and 	XG18345 	(g31224,g23932,g30280);
	or 	XG18346 	(g33321,g32182,g29712);
	or 	XG18347 	(g30515,g22036,g30223);
	nor 	XG18348 	(g33432,g6978,g31997);
	nor 	XG18349 	(g33098,g4616,g31997);
	or 	XG18350 	(g33022,g21750,g32306);
	or 	XG18351 	(g33315,g32175,g29665);
	or 	XG18352 	(g33014,g18499,g32305);
	not 	XG18353 	(I29939,g31667);
	or 	XG18354 	(g33031,g21841,g32315);
	or 	XG18355 	(g30563,g22134,g29347);
	or 	XG18356 	(g33032,g21842,g32326);
	or 	XG18357 	(g30472,g21943,g30186);
	or 	XG18358 	(g32349,g31275,g29840);
	or 	XG18359 	(g32358,g31297,g29866);
	or 	XG18360 	(g30463,g21934,g30140);
	or 	XG18361 	(g30418,g21802,g29751);
	or 	XG18362 	(g33057,g22019,g31968);
	or 	XG18363 	(g33058,g22020,g31976);
	nor 	XG18364 	(g33088,g7224,g31997);
	nor 	XG18365 	(g33093,g4601,g31997);
	or 	XG18366 	(g32372,g31314,g29884);
	or 	XG18367 	(g30419,g21803,g29759);
	or 	XG18368 	(g32996,g18377,g32256);
	nor 	XG18369 	(g33449,g31950,g10311);
	nor 	XG18370 	(g33439,g4633,g31950);
	or 	XG18371 	(g32368,g31310,g29881);
	or 	XG18372 	(g30410,g21769,g29857);
	or 	XG18373 	(g31897,g24322,g31237);
	nor 	XG18374 	(g33095,g7236,g31997);
	nor 	XG18375 	(g33096,g4608,g31997);
	or 	XG18376 	(g30476,g21947,g30229);
	or 	XG18377 	(g33063,g22066,g31988);
	or 	XG18378 	(g32351,g31281,g29851);
	or 	XG18379 	(g30396,g21755,g29856);
	or 	XG18380 	(g30464,g21935,g30152);
	and 	XG18381 	(g31225,g21012,g30276);
	or 	XG18382 	(g30533,g22079,g30203);
	or 	XG18383 	(g30426,g21810,g29785);
	or 	XG18384 	(g32367,g31309,g29880);
	or 	XG18385 	(g30550,g22121,g30226);
	or 	XG18386 	(g30467,g21938,g30185);
	or 	XG18387 	(g30460,g21931,g30207);
	or 	XG18388 	(g30437,g21846,g29876);
	or 	XG18389 	(g33017,g18510,g32292);
	or 	XG18390 	(g30527,g22073,g30192);
	or 	XG18391 	(g33003,g18429,g32323);
	or 	XG18392 	(g32386,g29949,g31488);
	or 	XG18393 	(g32992,g18351,g32242);
	or 	XG18394 	(g30454,g21863,g29909);
	or 	XG18395 	(g30503,g22024,g30243);
	or 	XG18396 	(g33024,g21752,g32324);
	or 	XG18397 	(g32380,g31467,g29907);
	or 	XG18398 	(g30479,g21950,g29320);
	or 	XG18399 	(g33033,g21843,g32333);
	or 	XG18400 	(g30520,g22041,g30272);
	or 	XG18401 	(g30561,g22132,g30284);
	or 	XG18402 	(g33314,g32174,g29663);
	nor 	XG18403 	(g31498,g29540,g9030);
	nor 	XG18404 	(g31506,g29540,g4793);
	nor 	XG18405 	(g31116,g29540,g7892);
	nor 	XG18406 	(g31068,g29540,g4801);
	or 	XG18407 	(g32375,g31324,g29896);
	or 	XG18408 	(g30535,g22081,g30225);
	or 	XG18409 	(g33059,g22021,g31987);
	or 	XG18410 	(g30491,g21987,g30178);
	or 	XG18411 	(g33313,g32171,g29649);
	or 	XG18412 	(g30406,g21765,g29783);
	nor 	XG18413 	(g33437,g10275,g31997);
	or 	XG18414 	(g32989,g18326,g32241);
	or 	XG18415 	(g30485,g21981,g30166);
	nor 	XG18416 	(g33094,g4639,g31950);
	or 	XG18417 	(g30425,g21809,g29770);
	or 	XG18418 	(g30525,g22071,g30266);
	or 	XG18419 	(g30442,g21851,g29797);
	or 	XG18420 	(g30422,g21806,g29795);
	or 	XG18421 	(g30482,g21978,g30230);
	or 	XG18422 	(g30542,g22088,g29337);
	or 	XG18423 	(g33010,g18473,g32301);
	or 	XG18424 	(g30559,g22130,g30269);
	or 	XG18425 	(g30394,g21753,g29805);
	or 	XG18426 	(g30448,g21857,g29809);
	or 	XG18427 	(g30508,g22029,g30199);
	or 	XG18428 	(g30423,g21807,g29887);
	or 	XG18429 	(g30407,g21766,g29794);
	nor 	XG18430 	(g31507,g29556,g9064);
	or 	XG18431 	(g32355,g31286,g29855);
	or 	XG18432 	(g30415,g21799,g29843);
	or 	XG18433 	(g30514,g22035,g30211);
	or 	XG18434 	(g33018,g18525,g32312);
	or 	XG18435 	(g30478,g21949,g30248);
	not 	XG18436 	(g33127,g31950);
	or 	XG18437 	(g31896,g24305,g31242);
	or 	XG18438 	(g32998,g18393,g32300);
	or 	XG18439 	(g30484,g21980,g30154);
	and 	XG18440 	(g31229,g23949,g30288);
	and 	XG18441 	(g31226,g25218,g30282);
	or 	XG18442 	(g30408,g21767,g29806);
	or 	XG18443 	(g33026,g21795,g32307);
	nor 	XG18444 	(g33084,g7655,g31978);
	or 	XG18445 	(g30428,g21812,g29807);
	or 	XG18446 	(g33064,g22067,g31993);
	or 	XG18447 	(g30433,g21817,g29899);
	or 	XG18448 	(g30461,g21932,g30219);
	or 	XG18449 	(g30443,g21852,g29808);
	or 	XG18450 	(g30431,g21815,g29875);
	or 	XG18451 	(g33050,g21930,g31974);
	nor 	XG18452 	(g31126,g29540,g7928);
	or 	XG18453 	(g30537,g22083,g30246);
	or 	XG18454 	(g30500,g21996,g29326);
	or 	XG18455 	(g30493,g21989,g30198);
	not 	XG18456 	(g33413,g31971);
	or 	XG18457 	(g33027,g21796,g32314);
	or 	XG18458 	(g30417,g21801,g29874);
	or 	XG18459 	(g30509,g22030,g30210);
	or 	XG18460 	(g30470,g21941,g30165);
	or 	XG18461 	(g30409,g21768,g29842);
	not 	XG18462 	(I28925,g29987);
	and 	XG18463 	(g28722,g20738,g27955);
	and 	XG18464 	(g33849,g20387,g33262);
	and 	XG18465 	(g33647,g18878,g33390);
	and 	XG18466 	(g28660,g20623,g27824);
	and 	XG18467 	(g33844,g20327,g33257);
	and 	XG18468 	(g33640,g18831,g33387);
	and 	XG18469 	(g33883,g20589,g33294);
	and 	XG18470 	(g33879,g20566,g33289);
	and 	XG18471 	(g28327,g19785,g27365);
	and 	XG18472 	(g33871,g20546,g33281);
	and 	XG18473 	(g33848,g20384,g33261);
	and 	XG18474 	(g28683,g20649,g27876);
	and 	XG18475 	(g33106,g18990,g32408);
	and 	XG18476 	(g28639,g20597,g27767);
	and 	XG18477 	(g33881,g20586,g33292);
	and 	XG18478 	(g33865,g20526,g33275);
	and 	XG18479 	(g33101,g18976,g32398);
	and 	XG18480 	(g28343,g19799,g27380);
	and 	XG18481 	(g33840,g20267,g33253);
	and 	XG18482 	(g33858,g20448,g33268);
	and 	XG18483 	(g28703,g20680,g27925);
	and 	XG18484 	(g28360,g19861,g27401);
	and 	XG18485 	(g33882,g20587,g33293);
	and 	XG18486 	(g33870,g20545,g33280);
	and 	XG18487 	(g33847,g20383,g33260);
	and 	XG18488 	(g33885,g20609,g33296);
	and 	XG18489 	(g33646,g18876,g33389);
	nor 	XG18490 	(g33438,g4621,g31950);
	nor 	XG18491 	(g33448,g31950,g7785);
	nor 	XG18492 	(g31121,g29540,g4776);
	nor 	XG18493 	(g33090,g4593,g31997);
	nor 	XG18494 	(g33075,g7163,g31997);
	and 	XG18495 	(g30926,g21163,g29903);
	nor 	XG18496 	(g33092,g4332,g31978);
	and 	XG18497 	(g34523,g34351,g9162);
	and 	XG18498 	(g30920,g21024,g29889);
	nor 	XG18499 	(g31515,g29556,g4983);
	or 	XG18500 	(g32371,g31313,g29883);
	and 	XG18501 	(g30930,g23342,g29915);
	and 	XG18502 	(g30927,g24795,g29910);
	or 	XG18503 	(g33310,g32165,g29631);
	nor 	XG18504 	(g33109,g4584,g31997);
	not 	XG18505 	(g33804,g33250);
	and 	XG18506 	(g31219,g20875,g30265);
	and 	XG18507 	(g31182,g20682,g30240);
	and 	XG18508 	(g33311,g12925,g31942);
	and 	XG18509 	(g33305,g17811,g31935);
	and 	XG18510 	(g31230,g20751,g30285);
	and 	XG18511 	(g33269,g15582,g31970);
	and 	XG18512 	(g33264,g21306,g31965);
	or 	XG18513 	(g30495,g21991,g30222);
	or 	XG18514 	(g33012,g18483,g32274);
	or 	XG18515 	(g30453,g21862,g29902);
	or 	XG18516 	(g30496,g21992,g30231);
	or 	XG18517 	(g30439,g21848,g29761);
	or 	XG18518 	(g30519,g22040,g30264);
	or 	XG18519 	(g33007,g18455,g32331);
	or 	XG18520 	(g30505,g22026,g30168);
	or 	XG18521 	(g30546,g22117,g30277);
	or 	XG18522 	(g30548,g22119,g30204);
	or 	XG18523 	(g30403,g21762,g29750);
	or 	XG18524 	(g30558,g22129,g30258);
	or 	XG18525 	(g30475,g21946,g30220);
	or 	XG18526 	(g30429,g21813,g29844);
	or 	XG18527 	(g30549,g22120,g30215);
	or 	XG18528 	(g33013,g18484,g32283);
	or 	XG18529 	(g30451,g21860,g29877);
	or 	XG18530 	(g30488,g21984,g30197);
	or 	XG18531 	(g33004,g18431,g32246);
	or 	XG18532 	(g30416,g21800,g29858);
	or 	XG18533 	(g30545,g22116,g30268);
	or 	XG18534 	(g34438,g18150,g34348);
	or 	XG18535 	(g30552,g22123,g30283);
	or 	XG18536 	(g30517,g22038,g30244);
	or 	XG18537 	(g30529,g22075,g30212);
	or 	XG18538 	(g30486,g21982,g30177);
	or 	XG18539 	(g30497,g21993,g30242);
	and 	XG18540 	(g34524,g34359,g9083);
	nand 	XG18541 	(g34550,g12323,g34359,g626);
	or 	XG18542 	(g34537,g34084,g34324);
	nand 	XG18543 	(g34048,g7442,g10583,g33669);
	or 	XG18544 	(g30553,g22124,g30205);
	or 	XG18545 	(g30405,g21764,g29767);
	or 	XG18546 	(g30427,g21811,g29796);
	or 	XG18547 	(g30489,g21985,g30250);
	or 	XG18548 	(g30432,g21816,g29888);
	or 	XG18549 	(g33016,g18509,g32284);
	or 	XG18550 	(g30560,g22131,g30278);
	or 	XG18551 	(g30555,g22126,g30227);
	or 	XG18552 	(g30436,g21845,g29860);
	or 	XG18553 	(g30481,g21977,g30221);
	or 	XG18554 	(g30502,g22023,g30232);
	or 	XG18555 	(g30528,g22074,g30202);
	or 	XG18556 	(g33015,g18507,g32343);
	or 	XG18557 	(g30534,g22080,g30213);
	or 	XG18558 	(g30444,g21853,g29901);
	or 	XG18559 	(g30490,g21986,g30167);
	or 	XG18560 	(g33005,g18432,g32260);
	or 	XG18561 	(g33011,g18481,g32338);
	or 	XG18562 	(g30556,g22127,g30236);
	or 	XG18563 	(g30455,g21864,g30041);
	or 	XG18564 	(g30510,g22031,g30263);
	or 	XG18565 	(g30466,g21937,g30174);
	or 	XG18566 	(g33008,g18457,g32261);
	or 	XG18567 	(g30562,g22133,g30289);
	or 	XG18568 	(g30557,g22128,g30247);
	or 	XG18569 	(g30440,g21849,g29771);
	or 	XG18570 	(g30524,g22070,g30255);
	or 	XG18571 	(g30521,g22042,g29331);
	or 	XG18572 	(g30506,g22027,g30179);
	or 	XG18573 	(g30499,g21995,g30261);
	or 	XG18574 	(g30532,g22078,g30193);
	or 	XG18575 	(g30530,g22076,g30224);
	or 	XG18576 	(g30438,g21847,g29890);
	or 	XG18577 	(g30487,g21983,g30187);
	not 	XG18578 	(g34543,g34359);
	or 	XG18579 	(g30424,g21808,g29760);
	or 	XG18580 	(g30504,g22025,g30253);
	or 	XG18581 	(g30526,g22072,g30181);
	or 	XG18582 	(g30483,g21979,g30241);
	or 	XG18583 	(g30538,g22084,g30256);
	or 	XG18584 	(g34252,g18180,g34146);
	or 	XG18585 	(g30494,g21990,g30209);
	or 	XG18586 	(g32983,g18222,g31990);
	or 	XG18587 	(g30498,g21994,g30251);
	or 	XG18588 	(g30420,g21804,g29769);
	and 	XG18589 	(g34542,g20089,g34332);
	and 	XG18590 	(g34309,g34147,g13947);
	or 	XG18591 	(g34330,g33717,g34069);
	or 	XG18592 	(g34250,g21713,g34111);
	or 	XG18593 	(g34249,g21702,g34110);
	and 	XG18594 	(g34344,g20038,g34107);
	not 	XG18595 	(g34346,g34162);
	and 	XG18596 	(g34310,g34162,g14003);
	nor 	XG18597 	(g34354,g11083,g34162,g9003);
	or 	XG18598 	(g33039,g24312,g32187);
	not 	XG18599 	(g31578,I29199);
	nor 	XG18600 	(g33112,g32194,g31240);
	and 	XG18601 	(g33719,g19433,g33141);
	and 	XG18602 	(g33237,g25198,g32394);
	and 	XG18603 	(g33830,g20166,g33382);
	and 	XG18604 	(g33822,g20157,g33385);
	not 	XG18605 	(g30295,I28540);
	or 	XG18606 	(g33212,I30756,I30755,g32328);
	or 	XG18607 	(g33204,I30751,I30750,g32317);
	not 	XG18608 	(I27567,g28181);
	not 	XG18609 	(I27576,g28173);
	not 	XG18610 	(I28390,g29185);
	and 	XG18611 	(g33909,g10708,g33131);
	and 	XG18612 	(g33910,g7836,g33134);
	not 	XG18613 	(g32364,I29894);
	or 	XG18614 	(g33694,g33429,g32402);
	and 	XG18615 	(g33487,I31132,I31131,g32649);
	and 	XG18616 	(g33478,I31087,I31086,g32584);
	and 	XG18617 	(g33469,I31042,I31041,g32519);
	and 	XG18618 	(g33518,I31287,I31286,g32874);
	and 	XG18619 	(g33515,I31272,I31271,g32853);
	and 	XG18620 	(g33519,I31292,I31291,g32881);
	and 	XG18621 	(g33517,I31282,I31281,g32867);
	and 	XG18622 	(g33516,I31277,I31276,g32860);
	and 	XG18623 	(g33520,I31297,I31296,g32888);
	and 	XG18624 	(g33521,I31302,I31301,g32895);
	and 	XG18625 	(g33522,I31307,I31306,g32902);
	and 	XG18626 	(g33523,I31312,I31311,g32909);
	not 	XG18627 	(I27561,g28163);
	nand 	XG18628 	(g33838,g4369,g33083);
	not 	XG18629 	(g30072,I28301);
	not 	XG18630 	(g30569,I28838);
	not 	XG18631 	(I27579,g28184);
	not 	XG18632 	(g29368,I27730);
	or 	XG18633 	(g33197,I30746,I30745,g32342);
	or 	XG18634 	(g33219,I30761,I30760,g32335);
	and 	XG18635 	(g33528,I31337,I31336,g32946);
	and 	XG18636 	(g33506,I31227,I31226,g32788);
	and 	XG18637 	(g33507,I31232,I31231,g32795);
	and 	XG18638 	(g33500,I31197,I31196,g32744);
	and 	XG18639 	(g33502,I31207,I31206,g32758);
	and 	XG18640 	(g33509,I31242,I31241,g32809);
	and 	XG18641 	(g33513,I31262,I31261,g32837);
	and 	XG18642 	(g33527,I31332,I31331,g32939);
	and 	XG18643 	(g33512,I31257,I31256,g32830);
	and 	XG18644 	(g33510,I31247,I31246,g32816);
	and 	XG18645 	(g33511,I31252,I31251,g32823);
	and 	XG18646 	(g33524,I31317,I31316,g32918);
	and 	XG18647 	(g33531,I31352,I31351,g32967);
	and 	XG18648 	(g33530,I31347,I31346,g32960);
	and 	XG18649 	(g33499,I31192,I31191,g32737);
	and 	XG18650 	(g33503,I31212,I31211,g32765);
	and 	XG18651 	(g33498,I31187,I31186,g32730);
	and 	XG18652 	(g33508,I31237,I31236,g32802);
	and 	XG18653 	(g33525,I31322,I31321,g32925);
	and 	XG18654 	(g33497,I31182,I31181,g32723);
	and 	XG18655 	(g33526,I31327,I31326,g32932);
	and 	XG18656 	(g33504,I31217,I31216,g32772);
	and 	XG18657 	(g33501,I31202,I31201,g32751);
	and 	XG18658 	(g33529,I31342,I31341,g32953);
	and 	XG18659 	(g33489,I31142,I31141,g32665);
	and 	XG18660 	(g33493,I31162,I31161,g32693);
	and 	XG18661 	(g33492,I31157,I31156,g32686);
	and 	XG18662 	(g33491,I31152,I31151,g32679);
	and 	XG18663 	(g33490,I31147,I31146,g32672);
	and 	XG18664 	(g33495,I31172,I31171,g32707);
	and 	XG18665 	(g33488,I31137,I31136,g32658);
	and 	XG18666 	(g33494,I31167,I31166,g32700);
	and 	XG18667 	(g33484,I31117,I31116,g32628);
	and 	XG18668 	(g33486,I31127,I31126,g32642);
	and 	XG18669 	(g33485,I31122,I31121,g32635);
	and 	XG18670 	(g33479,I31092,I31091,g32593);
	and 	XG18671 	(g33481,I31102,I31101,g32607);
	and 	XG18672 	(g33482,I31107,I31106,g32614);
	and 	XG18673 	(g33480,I31097,I31096,g32600);
	and 	XG18674 	(g33496,I31177,I31176,g32714);
	and 	XG18675 	(g33461,I31002,I31001,g32463);
	and 	XG18676 	(g33464,I31017,I31016,g32484);
	and 	XG18677 	(g33463,I31012,I31011,g32477);
	and 	XG18678 	(g33462,I31007,I31006,g32470);
	and 	XG18679 	(g33466,I31027,I31026,g32498);
	and 	XG18680 	(g33468,I31037,I31036,g32512);
	and 	XG18681 	(g33467,I31032,I31031,g32505);
	and 	XG18682 	(g33475,I31072,I31071,g32563);
	and 	XG18683 	(g33471,I31052,I31051,g32535);
	and 	XG18684 	(g33477,I31082,I31081,g32577);
	and 	XG18685 	(g33476,I31077,I31076,g32570);
	and 	XG18686 	(g33470,I31047,I31046,g32528);
	and 	XG18687 	(g33473,I31062,I31061,g32549);
	and 	XG18688 	(g33472,I31057,I31056,g32542);
	not 	XG18689 	(g29371,I27735);
	not 	XG18690 	(g32383,I29913);
	not 	XG18691 	(I27549,g28161);
	or 	XG18692 	(g33709,g33441,g32414);
	nor 	XG18693 	(g33117,g32205,g31261);
	not 	XG18694 	(I27742,g28819);
	not 	XG18695 	(g32024,I29582);
	not 	XG18696 	(g29379,I27749);
	not 	XG18697 	(I29239,g29498);
	not 	XG18698 	(I29236,g29498);
	not 	XG18699 	(I27570,g28262);
	or 	XG18700 	(g33076,g32446,g32336);
	and 	XG18701 	(g33381,g32318,g11842);
	not 	XG18702 	(g30116,I28349);
	not 	XG18703 	(I27573,g28157);
	not 	XG18704 	(I29245,g29491);
	not 	XG18705 	(I29248,g29491);
	not 	XG18706 	(I27552,g28162);
	not 	XG18707 	(I27564,g28166);
	not 	XG18708 	(I27555,g28142);
	not 	XG18709 	(I28908,g30182);
	not 	XG18710 	(I27558,g28155);
	not 	XG18711 	(g33326,g32318);
	not 	XG18712 	(g32449,I29977);
	not 	XG18713 	(I27546,g29041);
	or 	XG18714 	(g33988,g18397,g33861);
	or 	XG18715 	(g34018,g18505,g33887);
	and 	XG18716 	(g33684,g13565,g33139);
	and 	XG18717 	(g33689,g11006,g33144);
	or 	XG18718 	(g32117,g30914,g24482);
	or 	XG18719 	(g33176,I30735,I30734,g32198);
	or 	XG18720 	(g33044,g24327,g32199);
	or 	XG18721 	(g33187,I30741,I30740,g32014);
	or 	XG18722 	(g33685,g33423,g32396);
	or 	XG18723 	(g33972,g18335,g33941);
	or 	XG18724 	(g32253,g31207,g24771);
	or 	XG18725 	(g32267,g31218,g31208);
	not 	XG18726 	(g33354,g32329);
	or 	XG18727 	(g33980,g18370,g33843);
	or 	XG18728 	(g33976,g18347,g33869);
	not 	XG18729 	(g32437,I29965);
	not 	XG18730 	(g33072,g31945);
	or 	XG18731 	(g33318,g32434,g31969);
	or 	XG18732 	(g33979,g18361,g33942);
	or 	XG18733 	(g33323,g32442,g31936);
	not 	XG18734 	(g32445,I29973);
	not 	XG18735 	(g33430,g32421);
	or 	XG18736 	(g34019,g18506,g33889);
	or 	XG18737 	(g33994,g18424,g33841);
	or 	XG18738 	(g34000,g18441,g33943);
	or 	XG18739 	(g33149,I30718,I30717,g32204);
	or 	XG18740 	(g33998,g18428,g33878);
	and 	XG18741 	(g33693,g13594,g33145);
	and 	XG18742 	(g33700,g11012,g33148);
	or 	XG18743 	(g34010,g18478,g33872);
	or 	XG18744 	(g33042,g24324,g32193);
	and 	XG18745 	(g33786,g20572,g33130);
	or 	XG18746 	(g33706,g33440,g32412);
	or 	XG18747 	(g33164,I30728,I30727,g32203);
	or 	XG18748 	(g33981,g18371,g33856);
	or 	XG18749 	(g34011,g18479,g33884);
	or 	XG18750 	(g34009,g18477,g33863);
	or 	XG18751 	(g33714,g33450,g32419);
	or 	XG18752 	(g33703,g33434,g32410);
	or 	XG18753 	(g34017,g18504,g33880);
	or 	XG18754 	(g34012,g18480,g33886);
	or 	XG18755 	(g31783,I29352,I29351);
	or 	XG18756 	(g33969,g18321,g33864);
	or 	XG18757 	(g33692,g33428,g32400);
	or 	XG18758 	(g33699,g33433,g32409);
	not 	XG18759 	(g30606,I28866);
	not 	XG18760 	(g32021,I29579);
	and 	XG18761 	(g33795,g20782,g33138);
	or 	XG18762 	(g33986,g18387,g33639);
	or 	XG18763 	(g33041,g24323,g32189);
	not 	XG18764 	(I28883,g30105);
	and 	XG18765 	(g33758,g20269,g33133);
	or 	XG18766 	(g33968,g18320,g33855);
	and 	XG18767 	(g33734,I31593,g33136,g7806);
	or 	XG18768 	(g34021,g18519,g33652);
	not 	XG18769 	(I29909,g31791);
	and 	XG18770 	(g33676,g7970,g33125);
	and 	XG18771 	(g33680,g4688,g33128);
	or 	XG18772 	(g34003,g18452,g33866);
	or 	XG18773 	(g33036,g24309,g32168);
	nand 	XG18774 	(g33394,g32426,g4474,g10159);
	or 	XG18775 	(g33970,g18322,g33868);
	and 	XG18776 	(g33532,I31357,I31356,g32974);
	and 	XG18777 	(g33505,I31222,I31221,g32779);
	and 	XG18778 	(g33514,I31267,I31266,g32844);
	and 	XG18779 	(g33474,I31067,I31066,g32556);
	and 	XG18780 	(g33465,I31022,I31021,g32491);
	and 	XG18781 	(g33483,I31112,I31111,g32621);
	or 	XG18782 	(g33983,g18373,g33877);
	or 	XG18783 	(g33040,g24313,g32164);
	or 	XG18784 	(g33038,g24311,g32184);
	or 	XG18785 	(g33037,g24310,g32177);
	or 	XG18786 	(g33966,g18318,g33837);
	or 	XG18787 	(g33043,g24325,g32195);
	or 	XG18788 	(g33996,g18426,g33862);
	or 	XG18789 	(g33975,g18346,g33860);
	or 	XG18790 	(g34002,g18451,g33857);
	or 	XG18791 	(g34016,g18503,g33867);
	or 	XG18792 	(g33045,g24328,g32206);
	or 	XG18793 	(g33974,g18345,g33846);
	or 	XG18794 	(g33967,g18319,g33842);
	or 	XG18795 	(g33977,g18348,g33876);
	or 	XG18796 	(g32132,g31479,g31487);
	or 	XG18797 	(g31591,g29353,g29358);
	not 	XG18798 	(g33375,g32377);
	not 	XG18799 	(g32433,I29961);
	and 	XG18800 	(g33421,g21455,g32374);
	and 	XG18801 	(g33412,g21411,g32362);
	and 	XG18802 	(g33901,g20920,g33317);
	and 	XG18803 	(g33087,g18888,g32391);
	and 	XG18804 	(g33722,g19445,g33175);
	and 	XG18805 	(g33721,g19440,g33163);
	and 	XG18806 	(g33406,g21399,g32355);
	and 	XG18807 	(g33411,g21410,g32361);
	and 	XG18808 	(g33416,g21423,g32370);
	and 	XG18809 	(g33897,g20777,g33315);
	and 	XG18810 	(g33082,g18877,g32389);
	and 	XG18811 	(g33405,g21398,g32354);
	and 	XG18812 	(g33074,g18830,g32387);
	and 	XG18813 	(g33410,g21409,g32360);
	and 	XG18814 	(g33401,g21381,g32349);
	and 	XG18815 	(g33893,g20706,g33313);
	and 	XG18816 	(g33263,g25481,g32393);
	and 	XG18817 	(g33927,g21412,g33094);
	and 	XG18818 	(g33718,g19432,g33147);
	and 	XG18819 	(g33720,g19439,g33161);
	and 	XG18820 	(g33715,g19416,g33135);
	and 	XG18821 	(g33408,g21407,g32358);
	and 	XG18822 	(g33414,g21421,g32367);
	and 	XG18823 	(g33081,g18875,g32388);
	and 	XG18824 	(g33896,g20771,g33314);
	and 	XG18825 	(g33404,g21397,g32353);
	and 	XG18826 	(g33402,g21395,g32351);
	and 	XG18827 	(g33392,g21362,g32344);
	and 	XG18828 	(g33446,g21607,g32385);
	and 	XG18829 	(g33399,g21379,g32346);
	and 	XG18830 	(g33407,g21406,g32357);
	and 	XG18831 	(g33073,g18828,g32386);
	and 	XG18832 	(g33892,g20701,g33312);
	and 	XG18833 	(g33403,g21396,g32352);
	and 	XG18834 	(g33400,g21380,g32347);
	and 	XG18835 	(g33418,g21425,g32372);
	and 	XG18836 	(g33425,g21466,g32380);
	and 	XG18837 	(g33091,g18897,g32392);
	and 	XG18838 	(g33904,g21059,g33321);
	and 	XG18839 	(g33422,g21456,g32375);
	and 	XG18840 	(g33900,g20913,g33316);
	and 	XG18841 	(g33420,g21454,g32373);
	and 	XG18842 	(g33086,g18887,g32390);
	and 	XG18843 	(g33415,g21422,g32368);
	and 	XG18844 	(g33409,g21408,g32359);
	not 	XG18845 	(g30991,I28925);
	and 	XG18846 	(g33730,g4633,g33127,g4621,g7202);
	and 	XG18847 	(g32029,g16482,g31318);
	and 	XG18848 	(g32031,g13464,g31372);
	and 	XG18849 	(g33832,g27991,g33088);
	and 	XG18850 	(g33833,g25852,g33093);
	or 	XG18851 	(g31288,g29914,g2955);
	and 	XG18852 	(g33911,g10725,g33137);
	and 	XG18853 	(g33915,g7846,g33140);
	and 	XG18854 	(g33687,g4878,g33132);
	and 	XG18855 	(g33681,g7991,g33129);
	or 	XG18856 	(g32288,g31229,g31226);
	or 	XG18857 	(g32280,g31225,g24790);
	and 	XG18858 	(g33742,I31600,g33142,g7828);
	and 	XG18859 	(g32032,g16515,g31373);
	and 	XG18860 	(g32036,g13486,g31469);
	and 	XG18861 	(g32403,g15842,g31117);
	and 	XG18862 	(g32411,g13469,g31119);
	and 	XG18863 	(g33111,g32421,g24005);
	and 	XG18864 	(g33810,g12768,g33427);
	and 	XG18865 	(g33802,g14545,g33097);
	and 	XG18866 	(g33690,g16280,g33146);
	and 	XG18867 	(g33697,g13330,g33160);
	and 	XG18868 	(g33114,g31945,g22139);
	and 	XG18869 	(g33809,g30184,g33432);
	and 	XG18870 	(g33814,g28144,g33098);
	and 	XG18871 	(g33790,g20643,g33108);
	and 	XG18872 	(g33787,g20595,g33103);
	and 	XG18873 	(g33760,g20328,g33143);
	not 	XG18874 	(g32407,I29939);
	or 	XG18875 	(g32279,g31224,g31220);
	and 	XG18876 	(g33784,g20531,g33107);
	or 	XG18877 	(g32252,g31206,g31183);
	and 	XG18878 	(g32428,g16261,g31133);
	and 	XG18879 	(g32420,g19533,g31127);
	and 	XG18880 	(g33902,g13202,g33085);
	and 	XG18881 	(g33898,g15655,g33419);
	nor 	XG18882 	(g34067,g11772,g33859);
	or 	XG18883 	(g32294,g31232,g31231);
	and 	XG18884 	(g33701,g16305,g33162);
	and 	XG18885 	(g33707,g13346,g33174);
	and 	XG18886 	(g33785,g20550,g33100);
	or 	XG18887 	(g32130,g30925,g30921);
	or 	XG18888 	(g32123,g30919,g30915);
	or 	XG18889 	(g33984,g18374,g33881);
	and 	XG18890 	(g33811,g17573,g33439);
	and 	XG18891 	(g33815,g12911,g33449);
	and 	XG18892 	(g33903,g19146,g33447);
	and 	XG18893 	(g33905,g15574,g33089);
	or 	XG18894 	(g32124,g30920,g24488);
	or 	XG18895 	(g33973,g18344,g33840);
	or 	XG18896 	(g34005,g18454,g33883);
	or 	XG18897 	(g33995,g18425,g33848);
	or 	XG18898 	(g29291,g18767,g28660);
	and 	XG18899 	(g32044,g20085,g31483);
	and 	XG18900 	(g32045,g16187,g31491);
	or 	XG18901 	(g33891,g33269,g33264);
	or 	XG18902 	(g33997,g18427,g33871);
	and 	XG18903 	(g33908,g18935,g33092);
	and 	XG18904 	(g33906,g22311,g33084);
	and 	XG18905 	(g32052,g13885,g31507);
	and 	XG18906 	(g32068,g10862,g31515);
	or 	XG18907 	(g33982,g18372,g33865);
	or 	XG18908 	(g32289,g31230,g24796);
	or 	XG18909 	(g33991,g18400,g33885);
	and 	XG18910 	(g32039,g20070,g31476);
	and 	XG18911 	(g32043,g16173,g31482);
	or 	XG18912 	(g29274,g18642,g28360);
	or 	XG18913 	(g33914,g33311,g33305);
	and 	XG18914 	(g33835,g33413,g4340);
	and 	XG18915 	(g33801,g25327,g33437);
	and 	XG18916 	(g33808,g22161,g33109);
	or 	XG18917 	(g32240,g31182,g24757);
	or 	XG18918 	(g32268,g31219,g24785);
	or 	XG18919 	(g33990,g18399,g33882);
	or 	XG18920 	(g34015,g18502,g33858);
	and 	XG18921 	(g33834,g29172,g33095);
	and 	XG18922 	(g33836,g27020,g33096);
	or 	XG18923 	(g29309,g18818,g28722);
	or 	XG18924 	(g29262,g18608,g28327);
	or 	XG18925 	(g33989,g18398,g33870);
	or 	XG18926 	(g34007,g18467,g33640);
	and 	XG18927 	(g32048,g13869,g31498);
	and 	XG18928 	(g32051,g10831,g31506);
	or 	XG18929 	(g29268,g18625,g28343);
	or 	XG18930 	(g29303,g18801,g28703);
	or 	XG18931 	(g34004,g18453,g33879);
	and 	XG18932 	(g32401,g13432,g31116);
	and 	XG18933 	(g32397,g15830,g31068);
	or 	XG18934 	(g34014,g18493,g33647);
	and 	XG18935 	(g32418,g16239,g31126);
	and 	XG18936 	(g32413,g19518,g31121);
	and 	XG18937 	(g34169,g31227,g33804);
	or 	XG18938 	(g33541,g18223,g33101);
	and 	XG18939 	(g33828,g24411,g33090);
	and 	XG18940 	(g33820,g26830,g33075);
	and 	XG18941 	(g33922,g7202,g33448);
	and 	XG18942 	(g33919,g10795,g33438);
	or 	XG18943 	(g33543,g18281,g33106);
	or 	XG18944 	(g32131,g30926,g24495);
	or 	XG18945 	(g32144,g30930,g30927);
	or 	XG18946 	(g34008,g18476,g33849);
	or 	XG18947 	(g33987,g18396,g33847);
	or 	XG18948 	(g29297,g18784,g28683);
	or 	XG18949 	(g29285,g18750,g28639);
	or 	XG18950 	(g34695,g34322,g34523);
	or 	XG18951 	(g33993,g18413,g33646);
	or 	XG18952 	(g34001,g18450,g33844);
	and 	XG18953 	(g33417,g21424,g32371);
	and 	XG18954 	(g33890,g20659,g33310);
	and 	XG18955 	(g34702,g20208,g34537);
	and 	XG18956 	(g34364,g24366,g34048);
	and 	XG18957 	(g34685,g34550,g14164);
	not 	XG18958 	(g34698,g34550);
	and 	XG18959 	(g34687,g34543,g14181);
	or 	XG18960 	(g34599,g18149,g34542);
	and 	XG18961 	(g34538,g20054,g34330);
	or 	XG18962 	(g34535,g34073,g34309);
	and 	XG18963 	(g34513,g34346,g9003);
	or 	XG18964 	(g34439,g18181,g34344);
	nand 	XG18965 	(g34545,g34354,g794,g11679);
	and 	XG18966 	(g34506,g34354,g8833);
	not 	XG18967 	(g34539,g34354);
	and 	XG18968 	(g33807,g25452,g33112);
	not 	XG18969 	(I29891,g31578);
	and 	XG18970 	(g33913,g9104,g33204,g23088);
	and 	XG18971 	(g33907,g9104,g33219,g23088);
	or 	XG18972 	(g33616,g24314,g33237);
	not 	XG18973 	(I30995,g32449);
	not 	XG18974 	(g30928,I28908);
	not 	XG18975 	(g31666,I29248);
	not 	XG18976 	(I28582,g30116);
	or 	XG18977 	(g34034,g18713,g33719);
	not 	XG18978 	(I31724,g33076);
	not 	XG18979 	(I31727,g33076);
	not 	XG18980 	(g31657,I29239);
	not 	XG18981 	(I28594,g29379);
	not 	XG18982 	(I30641,g32024);
	not 	XG18983 	(I30644,g32024);
	not 	XG18984 	(g29374,I27742);
	not 	XG18985 	(I30861,g32383);
	not 	XG18986 	(I28591,g29371);
	or 	XG18987 	(I31844,g33477,g33476,g33475,g33474);
	or 	XG18988 	(I31843,g33473,g33472,g33471,g33470);
	or 	XG18989 	(I31838,g33464,g33463,g33462,g33461);
	or 	XG18990 	(I31848,g33482,g33481,g33480,g33479);
	or 	XG18991 	(I31849,g33486,g33485,g33484,g33483);
	or 	XG18992 	(I31854,g33495,g33494,g33493,g33492);
	or 	XG18993 	(I31853,g33491,g33490,g33489,g33488);
	or 	XG18994 	(I31874,g33531,g33530,g33529,g33528);
	or 	XG18995 	(I31859,g33504,g33503,g33502,g33501);
	or 	XG18996 	(I31873,g33527,g33526,g33525,g33524);
	or 	XG18997 	(I31858,g33500,g33499,g33498,g33497);
	or 	XG18998 	(I31863,g33509,g33508,g33507,g33506);
	or 	XG18999 	(I31864,g33513,g33512,g33511,g33510);
	not 	XG19000 	(I31616,g33219);
	not 	XG19001 	(I31782,g33219);
	not 	XG19002 	(I31545,g33219);
	not 	XG19003 	(I31459,g33219);
	not 	XG19004 	(I31528,g33219);
	not 	XG19005 	(I31659,g33219);
	not 	XG19006 	(I31770,g33197);
	not 	XG19007 	(I31561,g33197);
	not 	XG19008 	(I31786,g33197);
	not 	XG19009 	(I31569,g33197);
	not 	XG19010 	(I31486,g33197);
	not 	XG19011 	(I31625,g33197);
	not 	XG19012 	(I28588,g29368);
	not 	XG19013 	(I28872,g30072);
	not 	XG19014 	(g34208,g33838);
	or 	XG19015 	(g33963,g18124,g33830);
	or 	XG19016 	(I31869,g33522,g33521,g33520,g33519);
	or 	XG19017 	(I31868,g33518,g33517,g33516,g33515);
	or 	XG19018 	(g34055,g33910,g33909);
	or 	XG19019 	(g33962,g18123,g33822);
	not 	XG19020 	(g30155,I28390);
	not 	XG19021 	(I31622,g33204);
	not 	XG19022 	(I31642,g33204);
	not 	XG19023 	(I31482,g33204);
	not 	XG19024 	(I31564,g33204);
	not 	XG19025 	(I31550,g33204);
	not 	XG19026 	(I31776,g33204);
	not 	XG19027 	(I31539,g33212);
	not 	XG19028 	(I31555,g33212);
	not 	XG19029 	(I31650,g33212);
	not 	XG19030 	(I31779,g33212);
	not 	XG19031 	(I31474,g33212);
	not 	XG19032 	(I31619,g33212);
	not 	XG19033 	(I29233,g30295);
	and 	XG19034 	(g34082,g19554,g33709);
	and 	XG19035 	(g34079,g19532,g33703);
	and 	XG19036 	(g34076,g19519,g33694);
	and 	XG19037 	(g34083,g19573,g33714);
	and 	XG19038 	(g33360,g20869,g32253);
	and 	XG19039 	(g33365,g20994,g32267);
	and 	XG19040 	(g33239,g19902,g32117);
	and 	XG19041 	(g33796,g25267,g33117);
	and 	XG19042 	(g34075,g19517,g33692);
	and 	XG19043 	(g34081,g19552,g33706);
	and 	XG19044 	(g34078,g19531,g33699);
	and 	XG19045 	(g34074,g19498,g33685);
	and 	XG19046 	(g34113,g19744,g33734);
	and 	XG19047 	(g32028,g29339,g30569);
	and 	XG19048 	(g31995,g30569,g28274);
	and 	XG19049 	(g33379,g32364,g30984);
	not 	XG19050 	(I30983,g32433);
	and 	XG19051 	(g33431,g32377,g32364);
	not 	XG19052 	(I29981,g31591);
	not 	XG19053 	(g32415,g31591);
	not 	XG19054 	(g32450,g31591);
	not 	XG19055 	(I30980,g32132);
	not 	XG19056 	(g33346,g32132);
	not 	XG19057 	(g33451,g32132);
	or 	XG19058 	(g34148,g19656,g33758);
	or 	XG19059 	(g34172,g19914,g33795);
	nand 	XG19060 	(g33679,g10308,g10737,g33394);
	or 	XG19061 	(I31839,g33468,g33467,g33466,g33465);
	nand 	XG19062 	(g33925,g4467,g4462,g33394);
	or 	XG19063 	(g34090,g33680,g33676);
	not 	XG19064 	(g32381,I29909);
	not 	XG19065 	(g30729,I28883);
	not 	XG19066 	(I30959,g32021);
	not 	XG19067 	(I30962,g32021);
	not 	XG19068 	(I29936,g30606);
	not 	XG19069 	(I29571,g31783);
	not 	XG19070 	(I31701,g33164);
	not 	XG19071 	(I31686,g33164);
	not 	XG19072 	(I31810,g33164);
	not 	XG19073 	(I31504,g33164);
	not 	XG19074 	(I31607,g33164);
	not 	XG19075 	(I31800,g33164);
	not 	XG19076 	(I31581,g33164);
	or 	XG19077 	(g34101,g33700,g33693);
	not 	XG19078 	(I31610,g33149);
	not 	XG19079 	(I31823,g33149);
	not 	XG19080 	(I31672,g33149);
	not 	XG19081 	(I31586,g33149);
	not 	XG19082 	(I31807,g33149);
	not 	XG19083 	(I31814,g33149);
	not 	XG19084 	(I30992,g32445);
	not 	XG19085 	(I31817,g33323);
	not 	XG19086 	(I31820,g33323);
	not 	XG19087 	(I31463,g33318);
	not 	XG19088 	(I31466,g33318);
	not 	XG19089 	(I30986,g32437);
	not 	XG19090 	(I31791,g33354);
	not 	XG19091 	(I31515,g33187);
	not 	XG19092 	(g33686,g33187);
	not 	XG19093 	(I31523,g33187);
	not 	XG19094 	(g33695,g33187);
	not 	XG19095 	(I31597,g33187);
	not 	XG19096 	(I31497,g33187);
	not 	XG19097 	(I31604,g33176);
	not 	XG19098 	(I31500,g33176);
	not 	XG19099 	(I31803,g33176);
	not 	XG19100 	(I31796,g33176);
	not 	XG19101 	(I31694,g33176);
	or 	XG19102 	(g34099,g33689,g33684);
	and 	XG19103 	(g33678,g22319,g10710,g33149);
	and 	XG19104 	(g33704,g22319,g10710,g33176);
	and 	XG19105 	(g33674,g22319,g10710,g33164);
	and 	XG19106 	(g33728,g33187,g10851,g22626);
	and 	XG19107 	(g33725,g33176,g10851,g22626);
	and 	XG19108 	(g33711,g22332,g10727,g33176);
	and 	XG19109 	(g33675,g22332,g10727,g33164);
	and 	XG19110 	(g33683,g22332,g10727,g33149);
	and 	XG19111 	(g33812,g9104,g33187,g23088);
	and 	XG19112 	(g33819,g9104,g33176,g23088);
	and 	XG19113 	(g33831,g9104,g33149,g23088);
	and 	XG19114 	(g33921,g19200,g9104,g33187);
	or 	XG19115 	(g33552,g18343,g33400);
	or 	XG19116 	(g33575,g18420,g33086);
	or 	XG19117 	(g33617,g24326,g33263);
	or 	XG19118 	(g34168,g19784,g33787);
	or 	XG19119 	(g34006,g18462,g33897);
	and 	XG19120 	(g34370,g10554,g34067);
	or 	XG19121 	(g33560,g18369,g33404);
	or 	XG19122 	(g33599,g18500,g33087);
	or 	XG19123 	(g33578,g18433,g33410);
	or 	XG19124 	(g33546,g18327,g33402);
	or 	XG19125 	(g34167,g19768,g33786);
	or 	XG19126 	(g33545,g18324,g33399);
	or 	XG19127 	(g33551,g18342,g33446);
	or 	XG19128 	(g33999,g18436,g33893);
	or 	XG19129 	(g33584,g18449,g33406);
	or 	XG19130 	(g33586,g18459,g33416);
	or 	XG19131 	(g33561,g18376,g33408);
	or 	XG19132 	(g33544,g18317,g33392);
	or 	XG19133 	(g33992,g18408,g33900);
	or 	XG19134 	(g34103,g33707,g33701);
	nand 	XG19135 	(g33933,g12796,g12819,g12491,g33394);
	nand 	XG19136 	(g33930,g9848,g12767,g33394);
	or 	XG19137 	(g33585,g18456,g33411);
	or 	XG19138 	(g34170,g19855,g33790);
	or 	XG19139 	(g34013,g18488,g33901);
	or 	XG19140 	(g34231,g33902,g33898);
	or 	XG19141 	(g33119,g32428,g32420);
	or 	XG19142 	(g33600,g18501,g33418);
	or 	XG19143 	(g34026,g18682,g33715);
	not 	XG19144 	(I30901,g32407);
	or 	XG19145 	(g33583,g18448,g33074);
	or 	XG19146 	(g33562,g18379,g33414);
	or 	XG19147 	(g33607,g18526,g33091);
	or 	XG19148 	(g34028,g18684,g33720);
	or 	XG19149 	(g33570,g18405,g33420);
	or 	XG19150 	(g34193,g33814,g33809);
	or 	XG19151 	(g33577,g18430,g33405);
	or 	XG19152 	(g33985,g18382,g33896);
	or 	XG19153 	(g33601,g18508,g33422);
	or 	XG19154 	(g33553,g18350,g33403);
	or 	XG19155 	(g33568,g18395,g33409);
	or 	XG19156 	(g34020,g18514,g33904);
	or 	XG19157 	(g33554,g18353,g33407);
	or 	XG19158 	(g33592,g18475,g33412);
	or 	XG19159 	(g33569,g18402,g33415);
	or 	XG19160 	(g34100,g33697,g33690);
	or 	XG19161 	(g33602,g18511,g33425);
	or 	XG19162 	(g33576,g18423,g33401);
	or 	XG19163 	(g34025,g18672,g33927);
	or 	XG19164 	(g34190,g33810,g33802);
	or 	XG19165 	(g33559,g18368,g33073);
	or 	XG19166 	(g33594,g18485,g33421);
	or 	XG19167 	(g33116,g32411,g32403);
	or 	XG19168 	(g33231,g32036,g32032);
	or 	XG19169 	(g33591,g18474,g33082);
	or 	XG19170 	(g34036,g18715,g33722);
	or 	XG19171 	(g34035,g18714,g33721);
	or 	XG19172 	(g33567,g18394,g33081);
	or 	XG19173 	(g34027,g18683,g33718);
	or 	XG19174 	(g34095,g33687,g33681);
	or 	XG19175 	(g34057,g33915,g33911);
	or 	XG19176 	(g34204,g33833,g33832);
	or 	XG19177 	(g33227,g32031,g32029);
	or 	XG19178 	(g33978,g18356,g33892);
	not 	XG19179 	(g32438,g30991);
	not 	XG19180 	(g31937,g30991);
	not 	XG19181 	(I29969,g30991);
	and 	XG19182 	(g33374,g21221,g32289);
	and 	XG19183 	(g33376,g21268,g32294);
	and 	XG19184 	(g34117,g19755,g33742);
	and 	XG19185 	(g33242,g19931,g32123);
	and 	XG19186 	(g33366,g21010,g32268);
	and 	XG19187 	(g33370,g21139,g32279);
	and 	XG19188 	(g34226,g21467,g33914);
	and 	XG19189 	(g34211,g21349,g33891);
	and 	XG19190 	(g34066,g19352,g33730);
	and 	XG19191 	(g33359,g20853,g32252);
	and 	XG19192 	(g33353,g20732,g32240);
	and 	XG19193 	(g33243,g19947,g32124);
	and 	XG19194 	(g33247,g19980,g32130);
	and 	XG19195 	(g34774,g20180,g34695);
	and 	XG19196 	(g33371,g21155,g32280);
	and 	XG19197 	(g33373,g21205,g32288);
	and 	XG19198 	(g33249,g20026,g32144);
	and 	XG19199 	(g33248,g19996,g32131);
	or 	XG19200 	(g34166,g19752,g33785);
	or 	XG19201 	(g34149,g19674,g33760);
	or 	XG19202 	(g34158,g19740,g33784);
	or 	XG19203 	(g34064,g33922,g33919);
	or 	XG19204 	(g34199,g33828,g33820);
	not 	XG19205 	(I32352,g34169);
	or 	XG19206 	(g33118,g32418,g32413);
	or 	XG19207 	(g33115,g32401,g32397);
	or 	XG19208 	(g33238,g32051,g32048);
	or 	XG19209 	(g34206,g33836,g33834);
	or 	XG19210 	(g34189,g33808,g33801);
	or 	XG19211 	(g34207,g33304,g33835);
	or 	XG19212 	(g33234,g32043,g32039);
	or 	XG19213 	(g33240,g32068,g32052);
	or 	XG19214 	(g34046,g33908,g33906);
	or 	XG19215 	(g33236,g32045,g32044);
	or 	XG19216 	(g34043,g33905,g33903);
	or 	XG19217 	(g34194,g33815,g33811);
	or 	XG19218 	(g33593,g18482,g33417);
	or 	XG19219 	(g34440,g24226,g34364);
	or 	XG19220 	(g34724,g18152,g34702);
	or 	XG19221 	(g33971,g18330,g33890);
	and 	XG19222 	(g34742,g34698,g9000);
	or 	XG19223 	(g34762,g34524,g34687);
	or 	XG19224 	(g34600,g18182,g34538);
	and 	XG19225 	(g34700,g20129,g34535);
	or 	XG19226 	(g34693,g34310,g34513);
	not 	XG19227 	(g34697,g34545);
	and 	XG19228 	(g34684,g34545,g14178);
	nor 	XG19229 	(g34703,g11083,g34545,g8899);
	and 	XG19230 	(g34679,g34539,g14093);
	not 	XG19231 	(g32363,I29891);
	or 	XG19232 	(g34024,g24331,g33807);
	and 	XG19233 	(g34291,g19366,g34055);
	not 	XG19234 	(g31655,I29233);
	not 	XG19235 	(g33766,I31619);
	not 	XG19236 	(g33641,I31474);
	not 	XG19237 	(g33917,I31779);
	not 	XG19238 	(g33806,I31650);
	not 	XG19239 	(g33708,I31555);
	not 	XG19240 	(g33698,I31539);
	not 	XG19241 	(g33916,I31776);
	not 	XG19242 	(g33705,I31550);
	not 	XG19243 	(g33713,I31564);
	not 	XG19244 	(g33648,I31482);
	not 	XG19245 	(g33800,I31642);
	not 	XG19246 	(g33772,I31622);
	not 	XG19247 	(I28897,g30155);
	or 	XG19248 	(g33953,I31849,I31848,g33487);
	or 	XG19249 	(g33952,I31844,I31843,g33478);
	not 	XG19250 	(I32364,g34208);
	not 	XG19251 	(g30610,I28872);
	not 	XG19252 	(g33778,I31625);
	not 	XG19253 	(g33653,I31486);
	not 	XG19254 	(g33716,I31569);
	not 	XG19255 	(g33920,I31786);
	not 	XG19256 	(g33712,I31561);
	not 	XG19257 	(g33912,I31770);
	not 	XG19258 	(g33813,I31659);
	not 	XG19259 	(g33691,I31528);
	not 	XG19260 	(g33631,I31459);
	not 	XG19261 	(g33702,I31545);
	not 	XG19262 	(g33918,I31782);
	not 	XG19263 	(g33761,I31616);
	or 	XG19264 	(g33951,I31839,I31838,g33469);
	not 	XG19265 	(g33335,I30861);
	not 	XG19266 	(I28597,g29374);
	not 	XG19267 	(g33080,I30644);
	not 	XG19268 	(g32382,g31657);
	not 	XG19269 	(g33875,I31727);
	not 	XG19270 	(g32384,g31666);
	not 	XG19271 	(I29444,g30928);
	not 	XG19272 	(g33459,I30995);
	not 	XG19273 	(g34156,g33907);
	not 	XG19274 	(g34181,g33913);
	and 	XG19275 	(g34179,g24372,g33686);
	and 	XG19276 	(g34183,g24385,g33695);
	or 	XG19277 	(g33620,g18774,g33360);
	not 	XG19278 	(g33845,I31694);
	not 	XG19279 	(g33926,I31796);
	not 	XG19280 	(g33929,I31803);
	not 	XG19281 	(g33665,I31500);
	not 	XG19282 	(g33744,I31604);
	not 	XG19283 	(g33661,I31497);
	not 	XG19284 	(g33736,I31597);
	not 	XG19285 	(g33688,I31523);
	not 	XG19286 	(g33682,I31515);
	or 	XG19287 	(g33621,g18775,g33365);
	or 	XG19288 	(g34267,g18728,g34079);
	not 	XG19289 	(g33923,I31791);
	not 	XG19290 	(g33456,I30986);
	not 	XG19291 	(g33637,I31466);
	not 	XG19292 	(g33936,I31820);
	not 	XG19293 	(g33458,I30992);
	not 	XG19294 	(g33934,I31814);
	not 	XG19295 	(g33931,I31807);
	not 	XG19296 	(g33729,I31586);
	not 	XG19297 	(g33827,I31672);
	not 	XG19298 	(g33937,I31823);
	not 	XG19299 	(g33755,I31610);
	not 	XG19300 	(g33726,I31581);
	not 	XG19301 	(g33928,I31800);
	not 	XG19302 	(g33750,I31607);
	not 	XG19303 	(g33670,I31504);
	not 	XG19304 	(g33932,I31810);
	not 	XG19305 	(g33839,I31686);
	not 	XG19306 	(g33850,I31701);
	or 	XG19307 	(g34260,g18680,g34113);
	not 	XG19308 	(g32015,I29571);
	not 	XG19309 	(g32404,I29936);
	not 	XG19310 	(g33436,I30962);
	or 	XG19311 	(g33609,g18615,g33239);
	or 	XG19312 	(g34264,g18701,g34081);
	not 	XG19313 	(I29447,g30729);
	or 	XG19314 	(g34266,g18719,g34076);
	or 	XG19315 	(g34261,g18688,g34074);
	or 	XG19316 	(g34263,g18699,g34078);
	not 	XG19317 	(I30686,g32381);
	or 	XG19318 	(g34268,g18730,g34082);
	or 	XG19319 	(g33958,I31874,I31873,g33532);
	or 	XG19320 	(g33955,I31859,I31858,g33505);
	or 	XG19321 	(g33956,I31864,I31863,g33514);
	or 	XG19322 	(g33954,I31854,I31853,g33496);
	or 	XG19323 	(g34023,g24320,g33796);
	or 	XG19324 	(g33957,I31869,I31868,g33523);
	or 	XG19325 	(g34262,g18697,g34075);
	or 	XG19326 	(g34269,g18732,g34083);
	not 	XG19327 	(g33888,g33346);
	not 	XG19328 	(g33454,I30980);
	not 	XG19329 	(g33424,g32415);
	not 	XG19330 	(g32453,I29981);
	or 	XG19331 	(g33791,g32430,g33379);
	not 	XG19332 	(g33455,I30983);
	and 	XG19333 	(g33743,g19574,g33119);
	and 	XG19334 	(g33731,g19520,g33116);
	and 	XG19335 	(g33803,g20071,g33231);
	and 	XG19336 	(g34337,g19881,g34095);
	and 	XG19337 	(g34342,g19998,g34103);
	and 	XG19338 	(g34295,g19370,g34057);
	and 	XG19339 	(g34341,g19952,g34101);
	and 	XG19340 	(g34390,g21069,g34172);
	and 	XG19341 	(g34382,g20618,g34167);
	and 	XG19342 	(g34385,g20642,g34168);
	and 	XG19343 	(g34363,g20389,g34148);
	and 	XG19344 	(g34389,g20715,g34170);
	and 	XG19345 	(g34395,g21336,g34193);
	and 	XG19346 	(g34410,g21427,g34204);
	and 	XG19347 	(g34279,g19208,g34231);
	and 	XG19348 	(g34120,g25158,g33930);
	and 	XG19349 	(g34173,g24368,g33679);
	and 	XG19350 	(g34116,g25140,g33933);
	and 	XG19351 	(g34171,g24360,g33925);
	and 	XG19352 	(g34394,g21305,g34190);
	and 	XG19353 	(g33798,g20058,g33227);
	and 	XG19354 	(g34334,g19865,g34090);
	and 	XG19355 	(g34340,g19950,g34100);
	and 	XG19356 	(g34338,g19905,g34099);
	or 	XG19357 	(g33283,g30318,g31995);
	not 	XG19358 	(g32441,I29969);
	not 	XG19359 	(g33442,g31937);
	not 	XG19360 	(g33377,I30901);
	nor 	XG19361 	(g34496,g27648,g34370);
	not 	XG19362 	(g34192,g33921);
	not 	XG19363 	(g34132,g33831);
	not 	XG19364 	(g34124,g33819);
	not 	XG19365 	(g34197,g33812);
	not 	XG19366 	(g34053,g33683);
	not 	XG19367 	(g34044,g33675);
	not 	XG19368 	(g34062,g33711);
	not 	XG19369 	(g34070,g33725);
	not 	XG19370 	(g34068,g33728);
	not 	XG19371 	(g34042,g33674);
	not 	XG19372 	(g34060,g33704);
	not 	XG19373 	(g34049,g33678);
	or 	XG19374 	(g33610,g18616,g33242);
	or 	XG19375 	(g33612,g18633,g33247);
	or 	XG19376 	(g33618,g18757,g33353);
	or 	XG19377 	(g33624,g18808,g33371);
	or 	XG19378 	(g34258,g18675,g34211);
	or 	XG19379 	(g33627,g18826,g33376);
	or 	XG19380 	(g34257,g18674,g34226);
	or 	XG19381 	(g33619,g18758,g33359);
	or 	XG19382 	(g33623,g18792,g33370);
	or 	XG19383 	(g34790,g18151,g34774);
	or 	XG19384 	(g33622,g18791,g33366);
	or 	XG19385 	(g33626,g18825,g33374);
	or 	XG19386 	(g34259,g18679,g34066);
	not 	XG19387 	(g34345,I32352);
	or 	XG19388 	(g33613,g18649,g33248);
	or 	XG19389 	(g33614,g18650,g33249);
	or 	XG19390 	(g33625,g18809,g33373);
	or 	XG19391 	(g33611,g18632,g33243);
	or 	XG19392 	(g34265,g18711,g34117);
	and 	XG19393 	(g33829,g20164,g33240);
	and 	XG19394 	(g33818,g20113,g33236);
	and 	XG19395 	(g34380,g20571,g34158);
	and 	XG19396 	(g34381,g20594,g34166);
	and 	XG19397 	(g34365,g20451,g34149);
	and 	XG19398 	(g34401,g21383,g34199);
	and 	XG19399 	(g34393,g21304,g34189);
	and 	XG19400 	(g34281,g19276,g34043);
	and 	XG19401 	(g34414,g21457,g34206);
	and 	XG19402 	(g34284,g19351,g34046);
	and 	XG19403 	(g34396,g21337,g34194);
	and 	XG19404 	(g34415,g21458,g34207);
	and 	XG19405 	(g34301,g19415,g34064);
	and 	XG19406 	(g33735,g19553,g33118);
	and 	XG19407 	(g33821,g20153,g33238);
	and 	XG19408 	(g33727,g19499,g33115);
	and 	XG19409 	(g33816,g20096,g33234);
	or 	XG19410 	(g34826,g34685,g34742);
	and 	XG19411 	(g34842,g20168,g34762);
	or 	XG19412 	(g34725,g18183,g34700);
	and 	XG19413 	(g34771,g20147,g34693);
	and 	XG19414 	(g34741,g34697,g8899);
	or 	XG19415 	(g34761,g34506,g34679);
	and 	XG19416 	(g34743,g34703,g8951);
	not 	XG19417 	(g34766,g34703);
	not 	XG19418 	(I30766,g32363);
	and 	XG19419 	(g34109,g23708,g33918);
	and 	XG19420 	(g34097,g18957,g9104,g33772);
	and 	XG19421 	(g34102,g23599,g33912);
	and 	XG19422 	(g34112,g33778,g9104,g22957);
	and 	XG19423 	(g34096,g33772,g9104,g22957);
	and 	XG19424 	(g34087,g18957,g9104,g33766);
	and 	XG19425 	(g34086,g9104,g33766,g20114);
	and 	XG19426 	(g34106,g23675,g33917);
	and 	XG19427 	(g34063,g23121,g33806);
	and 	XG19428 	(g34212,g22689,g33761);
	and 	XG19429 	(g34214,g22689,g33772);
	and 	XG19430 	(g34216,g22689,g33778);
	and 	XG19431 	(g34213,g22689,g33766);
	and 	XG19432 	(g34050,g22942,g33772);
	and 	XG19433 	(g34045,g22942,g33766);
	and 	XG19434 	(g34054,g22942,g33778);
	and 	XG19435 	(g34230,g22942,g33761);
	and 	XG19436 	(g34215,g22670,g33778);
	and 	XG19437 	(g34061,g23076,g33800);
	and 	XG19438 	(g34104,g23639,g33916);
	and 	XG19439 	(g34085,g18957,g9104,g33761);
	and 	XG19440 	(g34108,g33766,g9104,g22957);
	and 	XG19441 	(g34091,g33761,g9104,g22957);
	and 	XG19442 	(g34065,g23148,g33813);
	and 	XG19443 	(g34114,g23742,g33920);
	and 	XG19444 	(g34105,g18957,g9104,g33778);
	and 	XG19445 	(g34186,g24396,g33705);
	and 	XG19446 	(g34178,g24361,g33712);
	and 	XG19447 	(g34184,g24388,g33698);
	and 	XG19448 	(g34182,g24384,g33691);
	and 	XG19449 	(g34180,g24373,g33716);
	and 	XG19450 	(g34187,g24397,g33708);
	and 	XG19451 	(g34191,g24404,g33713);
	and 	XG19452 	(g34185,g24389,g33702);
	not 	XG19453 	(g33391,g32384);
	not 	XG19454 	(g34188,g33875);
	not 	XG19455 	(g33388,g32382);
	not 	XG19456 	(g33658,g33080);
	nand 	XG19457 	(I31972,g33631,g33641);
	not 	XG19458 	(I32051,g33631);
	not 	XG19459 	(I32109,g33631);
	nand 	XG19460 	(I31983,g33648,g33653);
	not 	XG19461 	(I32106,g33653);
	not 	XG19462 	(I32062,g33653);
	not 	XG19463 	(I29438,g30610);
	not 	XG19464 	(g34358,I32364);
	or 	XG19465 	(g34461,g18681,g34291);
	not 	XG19466 	(g30917,I28897);
	not 	XG19467 	(g34094,g33772);
	not 	XG19468 	(I32059,g33648);
	not 	XG19469 	(I32119,g33648);
	not 	XG19470 	(I32056,g33641);
	not 	XG19471 	(I32096,g33641);
	not 	XG19472 	(I29585,g31655);
	not 	XG19473 	(I32158,g33791);
	not 	XG19474 	(I32161,g33791);
	and 	XG19475 	(g33071,g32404,g31591);
	not 	XG19476 	(I30998,g32453);
	and 	XG19477 	(g33110,g32415,g32404);
	and 	XG19478 	(g33899,g33335,g32132);
	not 	XG19479 	(I31829,g33454);
	and 	XG19480 	(g33924,g33346,g33335);
	or 	XG19481 	(g34402,g25084,g34179);
	or 	XG19482 	(g34405,g25103,g34183);
	and 	XG19483 	(g34319,g34156,g9535);
	not 	XG19484 	(g33120,I30686);
	not 	XG19485 	(g33635,g33436);
	not 	XG19486 	(I30971,g32015);
	nand 	XG19487 	(I32202,g33670,g33937);
	not 	XG19488 	(I32074,g33670);
	not 	XG19489 	(I32093,g33670);
	not 	XG19490 	(I32079,g33937);
	not 	XG19491 	(I32116,g33937);
	not 	XG19492 	(g34229,g33936);
	not 	XG19493 	(g34047,g33637);
	not 	XG19494 	(I32150,g33923);
	and 	XG19495 	(g34329,g34181,g14511);
	nand 	XG19496 	(I32185,g33661,g33665);
	not 	XG19497 	(I32067,g33661);
	not 	XG19498 	(I32103,g33661);
	not 	XG19499 	(I32089,g33665);
	not 	XG19500 	(I32071,g33665);
	and 	XG19501 	(g34196,g24485,g33682);
	and 	XG19502 	(g34203,g24537,g33726);
	and 	XG19503 	(g34205,g24541,g33729);
	and 	XG19504 	(g34198,g24491,g33688);
	and 	XG19505 	(g34080,g33750,g9104,g22957);
	and 	XG19506 	(g34093,g9104,g33755,g20114);
	and 	XG19507 	(g34072,g24872,g33839);
	and 	XG19508 	(g34119,g33755,g9104,g20516);
	and 	XG19509 	(g34092,g18957,g9104,g33750);
	and 	XG19510 	(g34115,g33750,g9104,g20516);
	and 	XG19511 	(g34138,g23828,g33929);
	and 	XG19512 	(g34141,g23828,g33932);
	and 	XG19513 	(g34143,g23828,g33934);
	and 	XG19514 	(g34217,g22876,g33736);
	and 	XG19515 	(g34223,g22876,g33744);
	and 	XG19516 	(g34228,g22942,g33750);
	and 	XG19517 	(g34225,g22942,g33744);
	and 	XG19518 	(g34219,g22942,g33736);
	and 	XG19519 	(g34224,g22670,g33736);
	and 	XG19520 	(g34218,g22670,g33744);
	and 	XG19521 	(g34098,g18957,g9104,g33744);
	and 	XG19522 	(g34139,g23314,g33827);
	and 	XG19523 	(g34089,g33744,g9104,g22957);
	and 	XG19524 	(g34088,g18957,g9104,g33736);
	and 	XG19525 	(g34077,g33736,g9104,g22957);
	and 	XG19526 	(g34136,g23293,g33850);
	and 	XG19527 	(g34133,g23958,g33845);
	and 	XG19528 	(g34135,g23802,g33926);
	and 	XG19529 	(g34140,g23802,g33931);
	and 	XG19530 	(g34137,g23802,g33928);
	or 	XG19531 	(g34253,g24300,g34171);
	and 	XG19532 	(g34706,g10570,g34496);
	or 	XG19533 	(g34463,g18686,g34338);
	or 	XG19534 	(g34465,g18712,g34295);
	or 	XG19535 	(g34467,g18717,g34341);
	or 	XG19536 	(g34254,g24301,g34116);
	or 	XG19537 	(g34468,g18718,g34342);
	or 	XG19538 	(g34037,g18734,g33803);
	or 	XG19539 	(g34039,g18736,g33743);
	or 	XG19540 	(g34444,g18546,g34389);
	not 	XG19541 	(I31535,g33377);
	or 	XG19542 	(g34255,g24302,g34120);
	or 	XG19543 	(g34456,g18669,g34395);
	or 	XG19544 	(g34462,g18685,g34334);
	or 	XG19545 	(g34449,g18662,g34279);
	or 	XG19546 	(g34464,g18687,g34340);
	or 	XG19547 	(g34256,g24303,g34173);
	or 	XG19548 	(g34443,g18545,g34385);
	or 	XG19549 	(g34447,g18552,g34363);
	or 	XG19550 	(g34445,g18548,g34382);
	or 	XG19551 	(g34446,g18550,g34390);
	or 	XG19552 	(g34038,g18735,g33731);
	or 	XG19553 	(g34466,g18716,g34337);
	or 	XG19554 	(g34453,g18666,g34410);
	or 	XG19555 	(g34029,g18703,g33798);
	or 	XG19556 	(g34457,g18670,g34394);
	not 	XG19557 	(I30989,g32441);
	not 	XG19558 	(I31491,g33283);
	not 	XG19559 	(I31494,g33283);
	and 	XG19560 	(g34397,g34068,g7673);
	and 	XG19561 	(g34367,g34042,g7404);
	and 	XG19562 	(g34388,g34062,g10802);
	and 	XG19563 	(g34298,g34132,g8679);
	and 	XG19564 	(g34371,g34044,g7450);
	not 	XG19565 	(I32639,g34345);
	and 	XG19566 	(g34386,g34060,g10800);
	and 	XG19567 	(g34398,g34070,g7684);
	and 	XG19568 	(g34335,g34197,g8461);
	and 	XG19569 	(g34287,g34124,g11370);
	and 	XG19570 	(g34333,g34192,g9984);
	and 	XG19571 	(g34378,g34053,g13095);
	and 	XG19572 	(g34375,g34049,g13077);
	or 	XG19573 	(g34458,g18671,g34396);
	or 	XG19574 	(g34450,g18663,g34281);
	or 	XG19575 	(g34441,g18540,g34381);
	or 	XG19576 	(g34040,g18737,g33818);
	or 	XG19577 	(g34033,g18708,g33821);
	or 	XG19578 	(g34041,g18739,g33829);
	or 	XG19579 	(g34448,g18553,g34365);
	or 	XG19580 	(g34455,g18668,g34284);
	or 	XG19581 	(g34442,g18542,g34380);
	or 	XG19582 	(g34032,g18706,g33816);
	or 	XG19583 	(g34454,g18667,g34414);
	or 	XG19584 	(g34030,g18704,g33727);
	or 	XG19585 	(g34031,g18705,g33735);
	or 	XG19586 	(g34452,g18665,g34401);
	or 	XG19587 	(g34460,g18677,g34301);
	or 	XG19588 	(g34459,g18673,g34415);
	or 	XG19589 	(g34451,g18664,g34393);
	and 	XG19590 	(g34867,g20145,g34826);
	or 	XG19591 	(g34849,g18154,g34842);
	or 	XG19592 	(g34791,g18184,g34771);
	or 	XG19593 	(g34819,g34684,g34741);
	and 	XG19594 	(g34841,g20080,g34761);
	and 	XG19595 	(g34811,g34766,g14165);
	not 	XG19596 	(g33228,I30766);
	or 	XG19597 	(g34300,g34230,g26864);
	or 	XG19598 	(g34352,g34109,g26079);
	not 	XG19599 	(g32027,I29585);
	or 	XG19600 	(g34278,g34212,g26829);
	not 	XG19601 	(g34145,I32096);
	not 	XG19602 	(g34121,I32056);
	nand 	XG19603 	(I31973,I31972,g33641);
	or 	XG19604 	(g34350,g34106,g26048);
	or 	XG19605 	(g34349,g34104,g26019);
	not 	XG19606 	(g34160,I32119);
	not 	XG19607 	(g34122,I32059);
	nand 	XG19608 	(I31985,I31983,g33648);
	not 	XG19609 	(I29441,g30917);
	or 	XG19610 	(g34321,g34065,g25866);
	or 	XG19611 	(g34399,g25067,g34178);
	or 	XG19612 	(g34347,g34102,g25986);
	or 	XG19613 	(g34314,g34061,g25831);
	or 	XG19614 	(g34280,g34213,g26833);
	or 	XG19615 	(g34407,g25124,g34185);
	not 	XG19616 	(I32607,g34358);
	or 	XG19617 	(g34353,g34114,g26088);
	not 	XG19618 	(g34123,I32062);
	not 	XG19619 	(g34151,I32106);
	not 	XG19620 	(g34152,I32109);
	not 	XG19621 	(g34118,I32051);
	nand 	XG19622 	(I31974,I31972,g33631);
	or 	XG19623 	(g34282,g34214,g26838);
	or 	XG19624 	(g34318,g34063,g25850);
	or 	XG19625 	(g34406,g25123,g34184);
	or 	XG19626 	(g34283,g34215,g26839);
	or 	XG19627 	(g34412,g25143,g34187);
	or 	XG19628 	(g34403,g25085,g34180);
	not 	XG19629 	(g34059,g33658);
	or 	XG19630 	(g34416,g25159,g34191);
	not 	XG19631 	(I31469,g33388);
	not 	XG19632 	(g34387,g34188);
	not 	XG19633 	(I31477,g33391);
	or 	XG19634 	(g34404,g25102,g34182);
	or 	XG19635 	(g34411,g25142,g34186);
	or 	XG19636 	(g34306,g34054,g25782);
	or 	XG19637 	(g34305,g34050,g25775);
	or 	XG19638 	(g34303,g34045,g25768);
	or 	XG19639 	(g34286,g34216,g26842);
	not 	XG19640 	(g34323,g34105);
	not 	XG19641 	(g34326,g34091);
	not 	XG19642 	(g34327,g34108);
	not 	XG19643 	(g34315,g34085);
	not 	XG19644 	(g34313,g34086);
	not 	XG19645 	(g34307,g34087);
	not 	XG19646 	(g34328,g34096);
	not 	XG19647 	(g34336,g34112);
	not 	XG19648 	(g34311,g34097);
	and 	XG19649 	(g34413,g22670,g34094);
	not 	XG19650 	(g34130,I32071);
	not 	XG19651 	(g34142,I32089);
	nand 	XG19652 	(I32186,I32185,g33665);
	not 	XG19653 	(g34150,I32103);
	not 	XG19654 	(g34126,I32067);
	nand 	XG19655 	(I32187,I32185,g33661);
	not 	XG19656 	(I32613,g34329);
	not 	XG19657 	(g34195,I32150);
	not 	XG19658 	(g34275,g34047);
	not 	XG19659 	(g34272,g34229);
	not 	XG19660 	(g34159,I32116);
	not 	XG19661 	(g34134,I32079);
	nand 	XG19662 	(I32203,I32202,g33937);
	not 	XG19663 	(g34144,I32093);
	not 	XG19664 	(g34131,I32074);
	nand 	XG19665 	(I32204,I32202,g33670);
	not 	XG19666 	(g33443,I30971);
	not 	XG19667 	(g34052,g33635);
	not 	XG19668 	(I31361,g33120);
	not 	XG19669 	(I32601,g34319);
	nand 	XG19670 	(I31984,I31983,g33653);
	or 	XG19671 	(g34153,g33451,g33899);
	not 	XG19672 	(g33944,I31829);
	or 	XG19673 	(g33628,g32450,g33071);
	not 	XG19674 	(g33460,I30998);
	not 	XG19675 	(g34202,I32161);
	and 	XG19676 	(g34482,g18917,g34405);
	and 	XG19677 	(g34478,g18904,g34402);
	not 	XG19678 	(g33660,I31494);
	not 	XG19679 	(g33457,I30989);
	or 	XG19680 	(g34294,g34225,g26855);
	or 	XG19681 	(g34376,g34140,g26301);
	or 	XG19682 	(g34331,g34072,g27121);
	or 	XG19683 	(g34368,g34135,g26274);
	or 	XG19684 	(g34273,g34203,g27765);
	or 	XG19685 	(g34274,g34205,g27822);
	not 	XG19686 	(g33696,I31535);
	or 	XG19687 	(g34289,g34218,g26847);
	or 	XG19688 	(g34372,g34137,g26287);
	or 	XG19689 	(g34421,g34198,g27686);
	or 	XG19690 	(g34369,g34136,g26279);
	or 	XG19691 	(g34288,g34217,g26846);
	or 	XG19692 	(g34293,g34224,g26854);
	or 	XG19693 	(g34374,g34139,g26294);
	or 	XG19694 	(g34373,g34138,g26292);
	or 	XG19695 	(g34290,g34219,g26848);
	or 	XG19696 	(g34417,g34196,g27678);
	or 	XG19697 	(g34377,g34141,g26304);
	or 	XG19698 	(g34292,g34223,g26853);
	or 	XG19699 	(g34379,g34143,g26312);
	or 	XG19700 	(g34366,g34133,g26257);
	nor 	XG19701 	(g34737,g30003,g34706);
	or 	XG19702 	(g34297,g34228,g26858);
	not 	XG19703 	(g34339,g34077);
	not 	XG19704 	(g34308,g34088);
	not 	XG19705 	(g34343,g34089);
	not 	XG19706 	(g34312,g34098);
	not 	XG19707 	(g34317,g34115);
	not 	XG19708 	(g34325,g34092);
	not 	XG19709 	(g34320,g34119);
	not 	XG19710 	(g34316,g34093);
	not 	XG19711 	(g34299,g34080);
	not 	XG19712 	(I32651,g34375);
	not 	XG19713 	(I32654,g34378);
	not 	XG19714 	(I32617,g34333);
	not 	XG19715 	(I32591,g34287);
	not 	XG19716 	(I32621,g34335);
	not 	XG19717 	(I32550,g34398);
	not 	XG19718 	(I32665,g34386);
	not 	XG19719 	(g34569,I32639);
	not 	XG19720 	(I32648,g34371);
	not 	XG19721 	(I32594,g34298);
	not 	XG19722 	(I32671,g34388);
	not 	XG19723 	(I32645,g34367);
	not 	XG19724 	(I32547,g34397);
	or 	XG19725 	(g34880,g18153,g34867);
	and 	XG19726 	(g34866,g20106,g34819);
	or 	XG19727 	(g34850,g18185,g34841);
	or 	XG19728 	(g34856,g34743,g34811);
	not 	XG19729 	(I31748,g33228);
	not 	XG19730 	(I31751,g33228);
	and 	XG19731 	(g34572,g33326,g34387);
	not 	XG19732 	(g33645,I31477);
	not 	XG19733 	(g33638,I31469);
	not 	XG19734 	(I32297,g34059);
	nand 	XG19735 	(g34051,I31974,I31973);
	not 	XG19736 	(I32222,g34118);
	not 	XG19737 	(g34420,g34152);
	nand 	XG19738 	(g34056,I31985,I31984);
	not 	XG19739 	(g34419,g34151);
	not 	XG19740 	(I32231,g34123);
	not 	XG19741 	(g34540,I32607);
	not 	XG19742 	(I32228,g34122);
	not 	XG19743 	(g34271,g34160);
	not 	XG19744 	(I32225,g34121);
	not 	XG19745 	(g34409,g34145);
	not 	XG19746 	(I30537,g32027);
	and 	XG19747 	(g34558,g20578,g34353);
	and 	XG19748 	(g34486,g18953,g34412);
	and 	XG19749 	(g34487,g18983,g34416);
	and 	XG19750 	(g34479,g18905,g34403);
	and 	XG19751 	(g34484,g18939,g34407);
	and 	XG19752 	(g34555,g20512,g34349);
	and 	XG19753 	(g34532,g19710,g34314);
	and 	XG19754 	(g34556,g20537,g34350);
	and 	XG19755 	(g34554,g20495,g34347);
	and 	XG19756 	(g34485,g18952,g34411);
	and 	XG19757 	(g34476,g18891,g34399);
	and 	XG19758 	(g34483,g18938,g34406);
	and 	XG19759 	(g34481,g18916,g34404);
	and 	XG19760 	(g34529,g19634,g34306);
	and 	XG19761 	(g34527,g19603,g34303);
	and 	XG19762 	(g34528,g19617,g34305);
	and 	XG19763 	(g34507,g19454,g34280);
	and 	XG19764 	(g34509,g19473,g34283);
	and 	XG19765 	(g34508,g19472,g34282);
	and 	XG19766 	(g34514,g19480,g34286);
	and 	XG19767 	(g34526,g19569,g34300);
	and 	XG19768 	(g34503,g19437,g34278);
	and 	XG19769 	(g34533,g19731,g34318);
	and 	XG19770 	(g34557,g20555,g34352);
	and 	XG19771 	(g34534,g19743,g34321);
	not 	XG19772 	(g34392,g34202);
	not 	XG19773 	(I32195,g33628);
	not 	XG19774 	(I32192,g33628);
	not 	XG19775 	(I32388,g34153);
	not 	XG19776 	(I32391,g34153);
	and 	XG19777 	(g33677,g31937,g33443);
	and 	XG19778 	(g33657,g33443,g30991);
	and 	XG19779 	(g34498,g34336,g13888);
	and 	XG19780 	(g34588,g34323,g26082);
	and 	XG19781 	(g34582,g34313,g7764);
	and 	XG19782 	(g34584,g34315,g24653);
	and 	XG19783 	(g34474,g34326,g20083);
	not 	XG19784 	(g34536,I32601);
	and 	XG19785 	(g34580,g34311,g29539);
	not 	XG19786 	(I32284,g34052);
	and 	XG19787 	(g34477,g34328,g26344);
	and 	XG19788 	(g34475,g34327,g27450);
	nand 	XG19789 	(g34227,I32204,I32203);
	not 	XG19790 	(I32240,g34131);
	not 	XG19791 	(g34408,g34144);
	not 	XG19792 	(I32243,g34134);
	not 	XG19793 	(g34270,g34159);
	and 	XG19794 	(g34492,g33430,g34272);
	or 	XG19795 	(g34494,g34413,g26849);
	and 	XG19796 	(g34577,g34307,g24577);
	not 	XG19797 	(I32274,g34195);
	not 	XG19798 	(g34544,I32613);
	nand 	XG19799 	(g34220,I32187,I32186);
	not 	XG19800 	(I32234,g34126);
	not 	XG19801 	(g34418,g34150);
	not 	XG19802 	(g34400,g34142);
	not 	XG19803 	(I32237,g34130);
	not 	XG19804 	(g34844,g34737);
	and 	XG19805 	(g34497,g33072,g34275);
	not 	XG19806 	(I31878,g33696);
	or 	XG19807 	(g34642,g18725,g34482);
	or 	XG19808 	(g34637,g18694,g34478);
	not 	XG19809 	(g34058,g33660);
	and 	XG19810 	(g34564,g17466,g34373);
	and 	XG19811 	(g34567,g17491,g34377);
	and 	XG19812 	(g34568,g17512,g34379);
	and 	XG19813 	(g34489,g19068,g34421);
	and 	XG19814 	(g34495,g19365,g34274);
	and 	XG19815 	(g34493,g19360,g34273);
	and 	XG19816 	(g34516,g19492,g34289);
	and 	XG19817 	(g34520,g19505,g34294);
	and 	XG19818 	(g34519,g19504,g34293);
	and 	XG19819 	(g34525,g19528,g34297);
	and 	XG19820 	(g34515,g19491,g34288);
	and 	XG19821 	(g34518,g19503,g34292);
	and 	XG19822 	(g34517,g19493,g34290);
	and 	XG19823 	(g34488,g18988,g34417);
	and 	XG19824 	(g34561,g17410,g34368);
	and 	XG19825 	(g34563,g17465,g34372);
	and 	XG19826 	(g34566,g17489,g34376);
	and 	XG19827 	(g34541,g20087,g34331);
	and 	XG19828 	(g34560,g17366,g34366);
	and 	XG19829 	(g34562,g17411,g34369);
	and 	XG19830 	(g34565,g17471,g34374);
	not 	XG19831 	(g34490,I32547);
	and 	XG19832 	(g34499,g34339,g31288);
	not 	XG19833 	(g34573,I32645);
	not 	XG19834 	(g34587,I32671);
	and 	XG19835 	(g34586,g34317,g11025);
	and 	XG19836 	(g34470,g34325,g7834);
	not 	XG19837 	(g34531,I32594);
	not 	XG19838 	(g34574,I32648);
	and 	XG19839 	(g34571,g34299,g27225);
	not 	XG19840 	(I32699,g34569);
	not 	XG19841 	(g34583,I32665);
	not 	XG19842 	(g34491,I32550);
	not 	XG19843 	(g34553,I32621);
	and 	XG19844 	(g34502,g34343,g26363);
	and 	XG19845 	(g34581,g34312,g22864);
	and 	XG19846 	(g34578,g34308,g24578);
	not 	XG19847 	(g34530,I32591);
	not 	XG19848 	(g34549,I32617);
	not 	XG19849 	(g34576,I32654);
	and 	XG19850 	(g34585,g34316,g24705);
	not 	XG19851 	(g34575,I32651);
	or 	XG19852 	(g34881,g18187,g34866);
	and 	XG19853 	(g34909,g20130,g34856);
	not 	XG19854 	(g33895,I31751);
	not 	XG19855 	(g34505,g34409);
	not 	XG19856 	(g34242,I32225);
	not 	XG19857 	(g34522,g34271);
	not 	XG19858 	(g34243,I32228);
	not 	XG19859 	(I32855,g34540);
	not 	XG19860 	(g34244,I32231);
	not 	XG19861 	(g34511,g34419);
	nand 	XG19862 	(I32431,g34051,g34056);
	not 	XG19863 	(g34512,g34420);
	not 	XG19864 	(g34241,I32222);
	not 	XG19865 	(g34296,I32297);
	not 	XG19866 	(I32170,g33638);
	or 	XG19867 	(g34708,g34572,g33381);
	not 	XG19868 	(I32173,g33645);
	not 	XG19869 	(g34246,I32237);
	not 	XG19870 	(g34501,g34400);
	or 	XG19871 	(g34619,g18581,g34528);
	not 	XG19872 	(g34510,g34418);
	not 	XG19873 	(g34245,I32234);
	nand 	XG19874 	(I32439,g34220,g34227);
	or 	XG19875 	(g34620,g18582,g34529);
	or 	XG19876 	(g34643,g18752,g34554);
	or 	XG19877 	(g34627,g18644,g34534);
	not 	XG19878 	(g34277,I32274);
	or 	XG19879 	(g34645,g18786,g34556);
	or 	XG19880 	(g34636,g18693,g34476);
	not 	XG19881 	(I32788,g34577);
	or 	XG19882 	(g34609,g18563,g34503);
	or 	XG19883 	(g34634,g18691,g34483);
	or 	XG19884 	(g34624,g18592,g34509);
	or 	XG19885 	(g34638,g18721,g34484);
	not 	XG19886 	(g34521,g34270);
	not 	XG19887 	(g34248,I32243);
	not 	XG19888 	(g34504,g34408);
	not 	XG19889 	(g34247,I32240);
	not 	XG19890 	(I32824,g34475);
	or 	XG19891 	(g34641,g18724,g34479);
	not 	XG19892 	(I32827,g34477);
	not 	XG19893 	(g34285,I32284);
	not 	XG19894 	(I32794,g34580);
	or 	XG19895 	(g34640,g18723,g34487);
	or 	XG19896 	(g34635,g18692,g34485);
	or 	XG19897 	(g34612,g18566,g34514);
	or 	XG19898 	(g34633,g18690,g34481);
	not 	XG19899 	(I32820,g34474);
	or 	XG19900 	(g34617,g18579,g34526);
	not 	XG19901 	(I32803,g34584);
	not 	XG19902 	(I32800,g34582);
	or 	XG19903 	(g34647,g18820,g34558);
	or 	XG19904 	(g34644,g18769,g34555);
	or 	XG19905 	(g34646,g18803,g34557);
	or 	XG19906 	(g34639,g18722,g34486);
	or 	XG19907 	(g34626,g18627,g34533);
	or 	XG19908 	(g34611,g18565,g34508);
	not 	XG19909 	(I32812,g34588);
	or 	XG19910 	(g34625,g18610,g34532);
	not 	XG19911 	(I32837,g34498);
	or 	XG19912 	(g34610,g18564,g34507);
	or 	XG19913 	(g34618,g18580,g34527);
	not 	XG19914 	(g34384,I32391);
	not 	XG19915 	(g34222,I32195);
	not 	XG19916 	(g34570,g34392);
	and 	XG19917 	(g34876,g20534,g34844);
	and 	XG19918 	(g34686,g19494,g34494);
	and 	XG19919 	(g34701,g20179,g34536);
	and 	XG19920 	(g34707,g20579,g34544);
	not 	XG19921 	(g34276,g34058);
	or 	XG19922 	(g34127,g32438,g33657);
	or 	XG19923 	(g34649,g34492,g33111);
	or 	XG19924 	(g34657,g34497,g33114);
	or 	XG19925 	(g34630,g15117,g34560);
	or 	XG19926 	(g34613,g18567,g34515);
	or 	XG19927 	(g34631,g15118,g34562);
	or 	XG19928 	(g34602,g18269,g34489);
	or 	XG19929 	(g34621,g18583,g34517);
	or 	XG19930 	(g34608,g15082,g34568);
	or 	XG19931 	(g34603,g15075,g34561);
	not 	XG19932 	(I32806,g34585);
	or 	XG19933 	(g34622,g18584,g34520);
	or 	XG19934 	(g34606,g15080,g34564);
	or 	XG19935 	(g34601,g18211,g34488);
	or 	XG19936 	(g34607,g15081,g34567);
	or 	XG19937 	(g34615,g18576,g34516);
	or 	XG19938 	(g34628,g18653,g34493);
	or 	XG19939 	(g34614,g18568,g34518);
	or 	XG19940 	(g34632,g15119,g34565);
	or 	XG19941 	(g34605,g15077,g34566);
	or 	XG19942 	(g34598,g18136,g34541);
	not 	XG19943 	(I32791,g34578);
	not 	XG19944 	(I32797,g34581);
	not 	XG19945 	(I32846,g34502);
	or 	XG19946 	(g34616,g18577,g34519);
	or 	XG19947 	(g34629,g18654,g34495);
	or 	XG19948 	(g34604,g15076,g34563);
	not 	XG19949 	(I32782,g34571);
	or 	XG19950 	(g34623,g18585,g34525);
	not 	XG19951 	(I32815,g34470);
	not 	XG19952 	(I32809,g34586);
	not 	XG19953 	(I32843,g34499);
	and 	XG19954 	(g34666,g19144,g34587);
	and 	XG19955 	(g34658,g18896,g34574);
	and 	XG19956 	(g34662,g18931,g34576);
	and 	XG19957 	(g34681,g19438,g34491);
	and 	XG19958 	(g34678,g19431,g34490);
	and 	XG19959 	(g34661,g18907,g34575);
	and 	XG19960 	(g34665,g19067,g34583);
	and 	XG19961 	(g34655,g18885,g34573);
	and 	XG19962 	(g34696,g20004,g34531);
	and 	XG19963 	(g34710,g20903,g34553);
	and 	XG19964 	(g34694,g19885,g34530);
	and 	XG19965 	(g34709,g17242,g34549);
	or 	XG19966 	(g34911,g18188,g34909);
	not 	XG19967 	(g34200,g33895);
	not 	XG19968 	(g34210,I32173);
	not 	XG19969 	(I32904,g34708);
	not 	XG19970 	(g34209,I32170);
	not 	XG19971 	(I32535,g34296);
	nand 	XG19972 	(I32433,I32431,g34051);
	not 	XG19973 	(I32452,g34241);
	not 	XG19974 	(I32775,g34512);
	not 	XG19975 	(I32763,g34511);
	not 	XG19976 	(I32461,g34244);
	not 	XG19977 	(g34699,I32855);
	not 	XG19978 	(I32458,g34243);
	not 	XG19979 	(I32766,g34522);
	not 	XG19980 	(I32455,g34242);
	not 	XG19981 	(I32770,g34505);
	not 	XG19982 	(g34423,g34222);
	not 	XG19983 	(g34559,g34384);
	not 	XG19984 	(g34689,I32837);
	not 	XG19985 	(g34676,I32812);
	not 	XG19986 	(g34672,I32800);
	not 	XG19987 	(g34673,I32803);
	nand 	XG19988 	(I32432,I32431,g34056);
	not 	XG19989 	(g34680,I32820);
	not 	XG19990 	(g34670,I32794);
	not 	XG19991 	(I32525,g34285);
	not 	XG19992 	(g34683,I32827);
	not 	XG19993 	(g34682,I32824);
	nand 	XG19994 	(I32440,I32439,g34227);
	not 	XG19995 	(I32470,g34247);
	not 	XG19996 	(I32874,g34504);
	not 	XG19997 	(I32473,g34248);
	not 	XG19998 	(I32871,g34521);
	not 	XG19999 	(g34668,I32788);
	not 	XG20000 	(I32476,g34277);
	not 	XG20001 	(I32464,g34245);
	not 	XG20002 	(I32752,g34510);
	not 	XG20003 	(I32878,g34501);
	not 	XG20004 	(I32467,g34246);
	nand 	XG20005 	(I32441,I32439,g34220);
	or 	XG20006 	(g34882,g18659,g34876);
	or 	XG20007 	(g34732,g18593,g34686);
	not 	XG20008 	(I32935,g34657);
	or 	XG20009 	(g34722,g18137,g34707);
	not 	XG20010 	(I32929,g34649);
	or 	XG20011 	(g34719,g18133,g34701);
	not 	XG20012 	(I32446,g34127);
	not 	XG20013 	(I32449,g34127);
	and 	XG20014 	(g34715,g33375,g34570);
	and 	XG20015 	(g34500,g30568,g34276);
	not 	XG20016 	(g34691,I32843);
	not 	XG20017 	(g34675,I32809);
	not 	XG20018 	(g34677,I32815);
	not 	XG20019 	(g34664,I32782);
	not 	XG20020 	(g34692,I32846);
	not 	XG20021 	(g34671,I32797);
	not 	XG20022 	(g34669,I32791);
	not 	XG20023 	(g34674,I32806);
	or 	XG20024 	(g34720,g18134,g34694);
	or 	XG20025 	(g34726,g18212,g34665);
	or 	XG20026 	(g34729,g18270,g34666);
	or 	XG20027 	(g34723,g18139,g34710);
	or 	XG20028 	(g34721,g18135,g34696);
	or 	XG20029 	(g34727,g18213,g34655);
	or 	XG20030 	(g34733,g18651,g34678);
	or 	XG20031 	(g34735,g15116,g34709);
	or 	XG20032 	(g34731,g18272,g34662);
	or 	XG20033 	(g34730,g18271,g34658);
	or 	XG20034 	(g34728,g18214,g34661);
	or 	XG20035 	(g34734,g18652,g34681);
	not 	XG20036 	(g34391,g34200);
	not 	XG20037 	(g34656,I32770);
	not 	XG20038 	(g34428,I32455);
	not 	XG20039 	(g34654,I32766);
	not 	XG20040 	(g34429,I32458);
	not 	XG20041 	(I32976,g34699);
	not 	XG20042 	(g34430,I32461);
	not 	XG20043 	(g34653,I32763);
	nand 	XG20044 	(g34422,I32433,I32432);
	not 	XG20045 	(g34659,I32775);
	not 	XG20046 	(g34427,I32452);
	not 	XG20047 	(g34480,I32535);
	not 	XG20048 	(I32305,g34209);
	not 	XG20049 	(g34736,I32904);
	not 	XG20050 	(I32309,g34210);
	not 	XG20051 	(g34432,I32467);
	not 	XG20052 	(g34716,I32878);
	not 	XG20053 	(g34648,I32752);
	not 	XG20054 	(g34431,I32464);
	nand 	XG20055 	(g34424,I32441,I32440);
	not 	XG20056 	(g34713,I32871);
	not 	XG20057 	(g34434,I32473);
	not 	XG20058 	(g34714,I32874);
	not 	XG20059 	(g34433,I32470);
	not 	XG20060 	(g34472,I32525);
	not 	XG20061 	(g34711,g34559);
	not 	XG20062 	(g34471,g34423);
	and 	XG20063 	(g34757,g19635,g34682);
	and 	XG20064 	(g34748,g19529,g34672);
	and 	XG20065 	(g34758,g19657,g34683);
	and 	XG20066 	(g34763,g19915,g34689);
	and 	XG20067 	(g34744,g19481,g34668);
	and 	XG20068 	(g34746,g19526,g34670);
	and 	XG20069 	(g34756,g19618,g34680);
	and 	XG20070 	(g34753,g19586,g34676);
	and 	XG20071 	(g34750,g19542,g34673);
	not 	XG20072 	(g34426,I32449);
	not 	XG20073 	(g34755,I32929);
	not 	XG20074 	(g34759,I32935);
	or 	XG20075 	(g34781,g34715,g33431);
	and 	XG20076 	(g34745,g19482,g34669);
	and 	XG20077 	(g34754,g19602,g34677);
	and 	XG20078 	(g34752,g19544,g34675);
	and 	XG20079 	(g34765,g20057,g34692);
	and 	XG20080 	(g34740,g19414,g34664);
	and 	XG20081 	(g34764,g20009,g34691);
	and 	XG20082 	(g34747,g19527,g34671);
	and 	XG20083 	(g34751,g19543,g34674);
	or 	XG20084 	(g34663,g34500,g32028);
	not 	XG20085 	(I32659,g34391);
	nand 	XG20086 	(I32516,g34422,g34424);
	not 	XG20087 	(g34304,I32309);
	not 	XG20088 	(I32985,g34736);
	not 	XG20089 	(g34302,I32305);
	not 	XG20090 	(I32840,g34480);
	not 	XG20091 	(I32675,g34427);
	not 	XG20092 	(I32947,g34659);
	not 	XG20093 	(I32960,g34653);
	not 	XG20094 	(I32684,g34430);
	not 	XG20095 	(g34778,I32976);
	not 	XG20096 	(I32681,g34429);
	not 	XG20097 	(I32956,g34654);
	not 	XG20098 	(I32678,g34428);
	not 	XG20099 	(I32953,g34656);
	and 	XG20100 	(g34667,g33424,g34471);
	and 	XG20101 	(g34782,g33888,g34711);
	not 	XG20102 	(I32834,g34472);
	not 	XG20103 	(I32693,g34433);
	not 	XG20104 	(I32973,g34714);
	not 	XG20105 	(I32696,g34434);
	not 	XG20106 	(I32950,g34713);
	not 	XG20107 	(I32687,g34431);
	not 	XG20108 	(I32967,g34648);
	not 	XG20109 	(I32970,g34716);
	not 	XG20110 	(I32690,g34432);
	or 	XG20111 	(g34801,g18588,g34756);
	or 	XG20112 	(g34792,g18569,g34750);
	or 	XG20113 	(g34794,g18571,g34746);
	or 	XG20114 	(g34803,g18590,g34758);
	or 	XG20115 	(g34806,g18595,g34763);
	or 	XG20116 	(g34795,g18572,g34753);
	not 	XG20117 	(I32991,g34759);
	or 	XG20118 	(g34802,g18589,g34757);
	or 	XG20119 	(g34793,g18570,g34744);
	not 	XG20120 	(I32988,g34755);
	or 	XG20121 	(g34805,g18594,g34748);
	not 	XG20122 	(g34473,g34426);
	not 	XG20123 	(I33020,g34781);
	or 	XG20124 	(g34799,g18578,g34751);
	or 	XG20125 	(g34797,g18574,g34747);
	or 	XG20126 	(g34798,g18575,g34754);
	or 	XG20127 	(g34804,g18591,g34740);
	or 	XG20128 	(g34800,g18586,g34752);
	or 	XG20129 	(g34796,g18573,g34745);
	or 	XG20130 	(g34807,g18596,g34764);
	or 	XG20131 	(g34808,g18599,g34765);
	not 	XG20132 	(I32938,g34663);
	not 	XG20133 	(g34579,I32659);
	not 	XG20134 	(g34769,I32953);
	not 	XG20135 	(g34590,I32678);
	not 	XG20136 	(g34770,I32956);
	not 	XG20137 	(g34591,I32681);
	not 	XG20138 	(I33053,g34778);
	not 	XG20139 	(I33056,g34778);
	not 	XG20140 	(g34592,I32684);
	not 	XG20141 	(g34772,I32960);
	nand 	XG20142 	(I32518,I32516,g34422);
	not 	XG20143 	(g34767,I32947);
	not 	XG20144 	(g34589,I32675);
	not 	XG20145 	(g34690,I32840);
	not 	XG20146 	(I32479,g34302);
	not 	XG20147 	(g34785,I32985);
	not 	XG20148 	(I32482,g34304);
	not 	XG20149 	(g34594,I32690);
	not 	XG20150 	(g34776,I32970);
	not 	XG20151 	(g34775,I32967);
	not 	XG20152 	(g34593,I32687);
	nand 	XG20153 	(I32517,I32516,g34424);
	not 	XG20154 	(g34768,I32950);
	not 	XG20155 	(g34596,I32696);
	not 	XG20156 	(g34777,I32973);
	not 	XG20157 	(g34595,I32693);
	not 	XG20158 	(g34688,I32834);
	or 	XG20159 	(g34843,g34782,g33924);
	or 	XG20160 	(g34783,g34667,g33110);
	not 	XG20161 	(g34660,g34473);
	not 	XG20162 	(g34786,I32988);
	not 	XG20163 	(g34787,I32991);
	not 	XG20164 	(g34810,I33020);
	not 	XG20165 	(g34760,I32938);
	not 	XG20166 	(I32868,g34579);
	nand 	XG20167 	(g34469,I32518,I32517);
	not 	XG20168 	(I32884,g34690);
	not 	XG20169 	(I33027,g34767);
	not 	XG20170 	(I33041,g34772);
	not 	XG20171 	(g34840,I33056);
	not 	XG20172 	(I33037,g34770);
	not 	XG20173 	(I33034,g34769);
	not 	XG20174 	(I33024,g34783);
	not 	XG20175 	(I33075,g34843);
	not 	XG20176 	(I32881,g34688);
	not 	XG20177 	(I33050,g34777);
	not 	XG20178 	(I33030,g34768);
	not 	XG20179 	(I33044,g34775);
	not 	XG20180 	(I33047,g34776);
	not 	XG20181 	(I33070,g34810);
	and 	XG20182 	(g34738,g33442,g34660);
	not 	XG20183 	(I32997,g34760);
	not 	XG20184 	(g34712,I32868);
	not 	XG20185 	(g34820,I33034);
	not 	XG20186 	(g34823,I33037);
	not 	XG20187 	(g34864,g34840);
	not 	XG20188 	(g34827,I33041);
	not 	XG20189 	(g34813,I33027);
	nand 	XG20190 	(I32756,g25779,g34469);
	not 	XG20191 	(g34718,I32884);
	not 	XG20192 	(g34833,I33047);
	not 	XG20193 	(g34830,I33044);
	not 	XG20194 	(g34816,I33030);
	not 	XG20195 	(g34836,I33050);
	not 	XG20196 	(g34717,I32881);
	not 	XG20197 	(g34851,I33075);
	not 	XG20198 	(g34812,I33024);
	not 	XG20199 	(g34848,I33070);
	not 	XG20200 	(g34789,I32997);
	or 	XG20201 	(g34809,g34738,g33677);
	not 	XG20202 	(I32909,g34712);
	nand 	XG20203 	(I32757,I32756,g34469);
	and 	XG20204 	(g34872,g19954,g34827);
	and 	XG20205 	(g34870,g19882,g34820);
	and 	XG20206 	(g34868,g19866,g34813);
	and 	XG20207 	(g34871,g19908,g34823);
	and 	XG20208 	(g34857,g34813,g16540);
	and 	XG20209 	(g34861,g34827,g16540);
	and 	XG20210 	(g34859,g34820,g16540);
	and 	XG20211 	(g34860,g34823,g16540);
	not 	XG20212 	(g34910,g34864);
	not 	XG20213 	(I33067,g34812);
	not 	XG20214 	(I33109,g34851);
	nand 	XG20215 	(I32758,I32756,g25779);
	and 	XG20216 	(g34862,g34830,g16540);
	and 	XG20217 	(g34863,g34833,g16540);
	and 	XG20218 	(g34858,g34816,g16540);
	and 	XG20219 	(g34865,g34836,g16540);
	and 	XG20220 	(g34874,g20060,g34833);
	and 	XG20221 	(g34873,g20046,g34830);
	and 	XG20222 	(g34869,g19869,g34816);
	and 	XG20223 	(g34875,g20073,g34836);
	not 	XG20224 	(I33079,g34809);
	not 	XG20225 	(g34739,I32909);
	not 	XG20226 	(I33182,g34910);
	nand 	XG20227 	(g34650,I32758,I32757);
	or 	XG20228 	(g34894,g21678,g34862);
	or 	XG20229 	(g34900,g21686,g34860);
	or 	XG20230 	(g34890,g21674,g34863);
	or 	XG20231 	(g34897,g21682,g34861);
	or 	XG20232 	(g34887,g21670,g34865);
	or 	XG20233 	(g34906,g21694,g34857);
	or 	XG20234 	(g34884,g21666,g34858);
	or 	XG20235 	(g34903,g21690,g34859);
	not 	XG20236 	(g34879,I33109);
	not 	XG20237 	(g34847,I33067);
	not 	XG20238 	(g34855,I33079);
	not 	XG20239 	(I32994,g34739);
	not 	XG20240 	(I32921,g34650);
	not 	XG20241 	(I32963,g34650);
	not 	XG20242 	(g34930,I33182);
	not 	XG20243 	(I33143,g34903);
	not 	XG20244 	(I33146,g34903);
	not 	XG20245 	(I33140,g34884);
	not 	XG20246 	(I33137,g34884);
	not 	XG20247 	(I33134,g34906);
	not 	XG20248 	(I33131,g34906);
	not 	XG20249 	(I33173,g34887);
	not 	XG20250 	(I33176,g34887);
	not 	XG20251 	(I33155,g34897);
	not 	XG20252 	(I33158,g34897);
	not 	XG20253 	(I33167,g34890);
	not 	XG20254 	(I33170,g34890);
	not 	XG20255 	(I33149,g34900);
	not 	XG20256 	(I33152,g34900);
	not 	XG20257 	(I33161,g34894);
	not 	XG20258 	(I33164,g34894);
	not 	XG20259 	(I33106,g34855);
	not 	XG20260 	(I33197,g34930);
	not 	XG20261 	(g34773,I32963);
	not 	XG20262 	(g34749,I32921);
	not 	XG20263 	(g34924,I33164);
	not 	XG20264 	(g34920,I33152);
	not 	XG20265 	(g34926,I33170);
	not 	XG20266 	(g34922,I33158);
	not 	XG20267 	(g34928,I33176);
	not 	XG20268 	(g34914,I33134);
	not 	XG20269 	(g34916,I33140);
	not 	XG20270 	(g34918,I33146);
	not 	XG20271 	(g34878,I33106);
	not 	XG20272 	(I32982,g34749);
	not 	XG20273 	(g34845,g34773);
	not 	XG20274 	(g34943,I33197);
	not 	XG20275 	(g34934,g34918);
	not 	XG20276 	(g34933,g34916);
	not 	XG20277 	(g34932,g34914);
	not 	XG20278 	(g34942,g34928);
	not 	XG20279 	(g34939,g34922);
	not 	XG20280 	(g34941,g34926);
	not 	XG20281 	(g34938,g34920);
	not 	XG20282 	(g34940,g34924);
	not 	XG20283 	(I33210,g34943);
	not 	XG20284 	(g34852,g34845);
	not 	XG20285 	(g34784,I32982);
	not 	XG20286 	(g34950,g34940);
	not 	XG20287 	(g34947,g34938);
	not 	XG20288 	(g34951,g34941);
	not 	XG20289 	(g34949,g34939);
	not 	XG20290 	(g34952,g34942);
	not 	XG20291 	(g34944,g34932);
	not 	XG20292 	(g34945,g34933);
	not 	XG20293 	(g34946,g34934);
	not 	XG20294 	(I33064,g34784);
	not 	XG20295 	(I33119,g34852);
	not 	XG20296 	(g34883,g34852);
	not 	XG20297 	(g34954,I33210);
	and 	XG20298 	(g34967,g23189,g34951);
	and 	XG20299 	(g34964,g23060,g34947);
	and 	XG20300 	(g34961,g23019,g34944);
	and 	XG20301 	(g34966,g23170,g34950);
	and 	XG20302 	(g34968,g23203,g34952);
	and 	XG20303 	(g34962,g23020,g34945);
	and 	XG20304 	(g34965,g23084,g34949);
	and 	XG20305 	(g34963,g23041,g34946);
	nor 	XG20306 	(g34912,g21370,g20242,g20277,g34883);
	not 	XG20307 	(I33214,g34954);
	not 	XG20308 	(g34893,I33119);
	not 	XG20309 	(g34846,I33064);
	or 	XG20310 	(g34977,g34966,g34873);
	or 	XG20311 	(g34970,g34961,g34868);
	or 	XG20312 	(g34975,g34964,g34871);
	or 	XG20313 	(g34978,g34967,g34874);
	or 	XG20314 	(g34979,g34968,g34875);
	or 	XG20315 	(g34971,g34962,g34869);
	or 	XG20316 	(g34976,g34965,g34872);
	or 	XG20317 	(g34974,g34963,g34870);
	not 	XG20318 	(I33103,g34846);
	not 	XG20319 	(I33179,g34893);
	or 	XG20320 	(g34931,g34912,g2984);
	not 	XG20321 	(I33264,g34978);
	not 	XG20322 	(I33255,g34975);
	not 	XG20323 	(I33246,g34970);
	not 	XG20324 	(I33261,g34977);
	not 	XG20325 	(I33252,g34974);
	not 	XG20326 	(I33258,g34976);
	not 	XG20327 	(I33249,g34971);
	not 	XG20328 	(I33267,g34979);
	not 	XG20329 	(g34929,I33179);
	not 	XG20330 	(g34877,I33103);
	and 	XG20331 	(g34955,g34320,g34931);
	not 	XG20332 	(g34987,I33261);
	not 	XG20333 	(g34982,I33246);
	not 	XG20334 	(g34985,I33255);
	not 	XG20335 	(g34988,I33264);
	not 	XG20336 	(g34989,I33267);
	not 	XG20337 	(g34983,I33249);
	not 	XG20338 	(g34986,I33258);
	not 	XG20339 	(g34984,I33252);
	not 	XG20340 	(I33189,g34929);
	not 	XG20341 	(I33285,g34988);
	not 	XG20342 	(I33276,g34985);
	not 	XG20343 	(I33270,g34982);
	not 	XG20344 	(I33282,g34987);
	not 	XG20345 	(I33218,g34955);
	not 	XG20346 	(I33273,g34984);
	not 	XG20347 	(I33279,g34986);
	not 	XG20348 	(I33291,g34983);
	not 	XG20349 	(I33288,g34989);
	not 	XG20350 	(g34935,I33189);
	not 	XG20351 	(g34960,I33218);
	not 	XG20352 	(g34994,I33282);
	not 	XG20353 	(g34990,I33270);
	not 	XG20354 	(g34992,I33276);
	not 	XG20355 	(g34995,I33285);
	not 	XG20356 	(g34996,I33288);
	not 	XG20357 	(g34997,I33291);
	not 	XG20358 	(g34993,I33279);
	not 	XG20359 	(g34991,I33273);
	and 	XG20360 	(g34953,g19957,g34935);
	and 	XG20361 	(g34948,g34935,g16540);
	and 	XG20362 	(g34969,g19570,g34960);
	or 	XG20363 	(g34957,g21662,g34948);
	or 	XG20364 	(g34980,g18587,g34969);
	not 	XG20365 	(I33235,g34957);
	not 	XG20366 	(I33232,g34957);
	not 	XG20367 	(g34973,I33235);
	not 	XG20368 	(g34981,g34973);
	not 	XG20369 	(g34998,g34981);
	and 	XG20370 	(g34999,g23085,g34998);
	or 	XG20371 	(g35000,g34999,g34953);
	not 	XG20372 	(I33297,g35000);
	not 	XG20373 	(g35001,I33297);
	not 	XG20374 	(I33300,g35001);
	not 	XG20375 	(g35002,I33300);
	not 	XG20376 	(g7243,I11892);
	not 	XG20377 	(g7245,I11896);
	not 	XG20378 	(g7257,I11903);
	not 	XG20379 	(g7260,I11908);
	not 	XG20380 	(g7540,I12026);
	not 	XG20381 	(g7916,I12300);
	not 	XG20382 	(g7946,I12314);
	not 	XG20383 	(g8132,I12411);
	not 	XG20384 	(g8178,I12437);
	not 	XG20385 	(g8215,I12451);
	not 	XG20386 	(g8235,I12463);
	not 	XG20387 	(g8277,I12483);
	not 	XG20388 	(g8279,I12487);
	not 	XG20389 	(g8283,I12493);
	not 	XG20390 	(g8291,I12503);
	not 	XG20391 	(g8342,I12519);
	not 	XG20392 	(g8344,I12523);
	not 	XG20393 	(g8353,I12530);
	not 	XG20394 	(g8358,I12541);
	not 	XG20395 	(g8398,I12563);
	not 	XG20396 	(g8403,I12568);
	not 	XG20397 	(g8416,I12580);
	not 	XG20398 	(g8475,I12608);
	not 	XG20399 	(g8719,I12719);
	not 	XG20400 	(g8783,I12761);
	not 	XG20401 	(g8784,I12764);
	not 	XG20402 	(g8785,I12767);
	not 	XG20403 	(g8786,I12770);
	not 	XG20404 	(g8787,I12773);
	not 	XG20405 	(g8788,I12776);
	not 	XG20406 	(g8789,I12779);
	not 	XG20407 	(g8839,I12819);
	not 	XG20408 	(g8870,I12837);
	not 	XG20409 	(g8915,I12884);
	not 	XG20410 	(g8916,I12887);
	not 	XG20411 	(g8917,I12890);
	not 	XG20412 	(g8918,I12893);
	not 	XG20413 	(g8919,I12896);
	not 	XG20414 	(g8920,I12899);
	not 	XG20415 	(g9019,I12950);
	not 	XG20416 	(g9048,I12963);
	not 	XG20417 	(g9251,I13037);
	not 	XG20418 	(g9497,I13166);
	not 	XG20419 	(g9553,I13202);
	not 	XG20420 	(g9555,I13206);
	not 	XG20421 	(g9615,I13236);
	not 	XG20422 	(g9617,I13240);
	not 	XG20423 	(g9680,I13276);
	not 	XG20424 	(g9682,I13280);
	not 	XG20425 	(g9741,I13317);
	not 	XG20426 	(g9743,I13321);
	not 	XG20427 	(g9817,I13374);
	not 	XG20428 	(g10122,I13623);
	not 	XG20429 	(g10306,I13726);
	not 	XG20430 	(g10500,I13875);
	not 	XG20431 	(g10527,I13892);
	not 	XG20432 	(g11349,I14365);
	not 	XG20433 	(g11388,I14395);
	not 	XG20434 	(g11418,I14424);
	not 	XG20435 	(g11447,I14450);
	not 	XG20436 	(g11678,I14563);
	not 	XG20437 	(g11770,I14619);
	not 	XG20438 	(g12184,I15036);
	not 	XG20439 	(g12238,I15102);
	not 	XG20440 	(g12300,I15144);
	not 	XG20441 	(g12350,I15190);
	not 	XG20442 	(g12368,I15208);
	not 	XG20443 	(g12422,I15238);
	not 	XG20444 	(g12470,I15284);
	or 	XG20445 	(g12832,g10348,g10347);
	not 	XG20446 	(g12919,I15536);
	not 	XG20447 	(g12923,I15542);
	not 	XG20448 	(g13039,I15663);
	not 	XG20449 	(g13049,I15677);
	not 	XG20450 	(g13068,I15697);
	not 	XG20451 	(g13085,I15717);
	not 	XG20452 	(g13099,I15732);
	not 	XG20453 	(g13259,I15824);
	not 	XG20454 	(g13272,I15837);
	not 	XG20455 	(g13865,I16168);
	not 	XG20456 	(g13881,I16181);
	not 	XG20457 	(g13895,I16193);
	not 	XG20458 	(g13906,I16201);
	not 	XG20459 	(g13926,I16217);
	not 	XG20460 	(g13966,I16246);
	not 	XG20461 	(g14096,I16328);
	not 	XG20462 	(g14125,I16345);
	not 	XG20463 	(g14147,I16357);
	not 	XG20464 	(g14167,I16371);
	not 	XG20465 	(g14189,I16391);
	not 	XG20466 	(g14201,I16401);
	not 	XG20467 	(g14217,I16417);
	not 	XG20468 	(g14421,I16575);
	not 	XG20469 	(g14451,I16606);
	not 	XG20470 	(g14518,I16639);
	not 	XG20471 	(g14597,I16713);
	not 	XG20472 	(g14635,I16741);
	not 	XG20473 	(g14662,I16762);
	not 	XG20474 	(g14673,I16770);
	not 	XG20475 	(g14694,I16795);
	not 	XG20476 	(g14705,I16803);
	not 	XG20477 	(g14738,I16821);
	not 	XG20478 	(g14749,I16829);
	not 	XG20479 	(g14779,I16847);
	not 	XG20480 	(g14828,I16875);
	not 	XG20481 	(g16603,I17787);
	not 	XG20482 	(g16624,I17814);
	not 	XG20483 	(g16627,I17819);
	not 	XG20484 	(g16656,I17852);
	not 	XG20485 	(g16659,I17857);
	not 	XG20486 	(g16686,I17892);
	not 	XG20487 	(g16693,I17901);
	not 	XG20488 	(g16718,I17932);
	not 	XG20489 	(g16722,I17938);
	not 	XG20490 	(g16744,I17964);
	not 	XG20491 	(g16748,I17970);
	not 	XG20492 	(g16775,I17999);
	not 	XG20493 	(g16874,I18066);
	not 	XG20494 	(g16924,I18092);
	not 	XG20495 	(g16955,I18107);
	not 	XG20496 	(g17291,I18276);
	not 	XG20497 	(g17316,I18293);
	not 	XG20498 	(g17320,I18297);
	not 	XG20499 	(g17400,I18333);
	not 	XG20500 	(g17404,I18337);
	not 	XG20501 	(g17423,I18360);
	not 	XG20502 	(g17519,I18460);
	not 	XG20503 	(g17577,I18504);
	not 	XG20504 	(g17580,I18509);
	not 	XG20505 	(g17604,I18555);
	not 	XG20506 	(g17607,I18560);
	not 	XG20507 	(g17639,I18600);
	not 	XG20508 	(g17646,I18609);
	not 	XG20509 	(g17649,I18614);
	not 	XG20510 	(g17674,I18647);
	not 	XG20511 	(g17678,I18653);
	not 	XG20512 	(g17685,I18662);
	not 	XG20513 	(g17688,I18667);
	not 	XG20514 	(g17711,I18694);
	not 	XG20515 	(g17715,I18700);
	not 	XG20516 	(g17722,I18709);
	not 	XG20517 	(g17739,I18728);
	not 	XG20518 	(g17743,I18734);
	not 	XG20519 	(g17760,I18752);
	not 	XG20520 	(g17764,I18758);
	not 	XG20521 	(g17778,I18778);
	not 	XG20522 	(g17787,I18795);
	not 	XG20523 	(g17813,I18813);
	not 	XG20524 	(g17819,I18825);
	not 	XG20525 	(g17845,I18835);
	not 	XG20526 	(g17871,I18845);
	not 	XG20527 	(g18092,I18882);
	not 	XG20528 	(g18094,I18888);
	not 	XG20529 	(g18095,I18891);
	not 	XG20530 	(g18096,I18894);
	not 	XG20531 	(g18097,I18897);
	not 	XG20532 	(g18098,I18900);
	not 	XG20533 	(g18099,I18903);
	not 	XG20534 	(g18100,I18906);
	not 	XG20535 	(g18101,I18909);
	not 	XG20536 	(g18881,I19671);
	not 	XG20537 	(g19334,I19818);
	not 	XG20538 	(g19357,I19837);
	not 	XG20539 	(g20049,I20318);
	not 	XG20540 	(g20557,I20647);
	not 	XG20541 	(g20652,I20744);
	not 	XG20542 	(g20654,I20750);
	not 	XG20543 	(g20763,I20816);
	not 	XG20544 	(g20899,I20861);
	not 	XG20545 	(g20901,I20867);
	not 	XG20546 	(g21176,I20954);
	not 	XG20547 	(g21245,I20982);
	not 	XG20548 	(g21270,I20999);
	not 	XG20549 	(g21292,I21033);
	not 	XG20550 	(g21698,g18562);
	not 	XG20551 	(g21727,I21300);
	not 	XG20552 	(g23002,I22177);
	not 	XG20553 	(g23190,I22286);
	not 	XG20554 	(g23612,I22745);
	not 	XG20555 	(g23652,I22785);
	not 	XG20556 	(g23683,I22816);
	not 	XG20557 	(g23759,I22886);
	or 	XG20558 	(g24151,g21661,g18088);
	not 	XG20559 	(g25114,I24278);
	not 	XG20560 	(g25167,I24331);
	not 	XG20561 	(g25219,I24393);
	not 	XG20562 	(g25259,I24445);
	or 	XG20563 	(g25582,g24152,g21662);
	or 	XG20564 	(g25583,g24153,g21666);
	or 	XG20565 	(g25584,g24154,g21670);
	or 	XG20566 	(g25585,g24155,g21674);
	or 	XG20567 	(g25586,g24156,g21678);
	or 	XG20568 	(g25587,g24157,g21682);
	or 	XG20569 	(g25588,g24158,g21686);
	or 	XG20570 	(g25589,g24159,g21690);
	or 	XG20571 	(g25590,g24160,g21694);
	not 	XG20572 	(g26801,I25511);
	or 	XG20573 	(g26875,g25575,g21652);
	or 	XG20574 	(g26876,g25576,g21655);
	or 	XG20575 	(g26877,g25577,g21658);
	not 	XG20576 	(g27831,I26406);
	or 	XG20577 	(g28030,g26874,g24018);
	or 	XG20578 	(g28041,g26878,g24145);
	or 	XG20579 	(g28042,g26879,g24148);
	not 	XG20580 	(g28753,I27235);
	not 	XG20581 	(g29210,I27546);
	not 	XG20582 	(g29211,I27549);
	not 	XG20583 	(g29212,I27552);
	not 	XG20584 	(g29213,I27555);
	not 	XG20585 	(g29214,I27558);
	not 	XG20586 	(g29215,I27561);
	not 	XG20587 	(g29216,I27564);
	not 	XG20588 	(g29217,I27567);
	not 	XG20589 	(g29218,I27570);
	not 	XG20590 	(g29219,I27573);
	not 	XG20591 	(g29220,I27576);
	not 	XG20592 	(g29221,I27579);
	not 	XG20593 	(g30327,I28582);
	not 	XG20594 	(g30329,I28588);
	not 	XG20595 	(g30330,I28591);
	not 	XG20596 	(g30331,I28594);
	not 	XG20597 	(g30332,I28597);
	not 	XG20598 	(g31521,I29182);
	not 	XG20599 	(g31656,I29236);
	not 	XG20600 	(g31665,I29245);
	or 	XG20601 	(g31793,g30317,g28031);
	not 	XG20602 	(g31860,I29438);
	not 	XG20603 	(g31861,I29441);
	not 	XG20604 	(g31862,I29444);
	not 	XG20605 	(g31863,I29447);
	not 	XG20606 	(g32185,I29717);
	or 	XG20607 	(g32429,g31794,g30318);
	or 	XG20608 	(g32454,g31795,g30322);
	not 	XG20609 	(g32975,I30537);
	not 	XG20610 	(g33079,I30641);
	not 	XG20611 	(g33435,I30959);
	not 	XG20612 	(g33533,I31361);
	not 	XG20613 	(g33636,I31463);
	not 	XG20614 	(g33659,I31491);
	not 	XG20615 	(g33874,I31724);
	not 	XG20616 	(g33894,I31748);
	not 	XG20617 	(g33935,I31817);
	or 	XG20618 	(g33945,g33455,g32430);
	or 	XG20619 	(g33946,g33456,g32434);
	or 	XG20620 	(g33947,g33457,g32438);
	or 	XG20621 	(g33948,g33458,g32442);
	or 	XG20622 	(g33949,g33459,g32446);
	or 	XG20623 	(g33950,g33460,g32450);
	not 	XG20624 	(g33959,I31878);
	not 	XG20625 	(g34201,I32158);
	not 	XG20626 	(g34221,I32192);
	or 	XG20627 	(g34232,g33944,g33451);
	or 	XG20628 	(g34233,g33951,g32455);
	or 	XG20629 	(g34234,g33952,g32520);
	or 	XG20630 	(g34235,g33953,g32585);
	or 	XG20631 	(g34236,g33954,g32650);
	or 	XG20632 	(g34237,g33955,g32715);
	or 	XG20633 	(g34238,g33956,g32780);
	or 	XG20634 	(g34239,g33957,g32845);
	or 	XG20635 	(g34240,g33958,g32910);
	not 	XG20636 	(g34383,I32388);
	not 	XG20637 	(g34425,I32446);
	not 	XG20638 	(g34435,I32476);
	not 	XG20639 	(g34436,I32479);
	not 	XG20640 	(g34437,I32482);
	not 	XG20641 	(g34597,I32699);
	not 	XG20642 	(g34788,I32994);
	not 	XG20643 	(g34839,I33053);
	not 	XG20644 	(g34913,I33131);
	not 	XG20645 	(g34915,I33137);
	not 	XG20646 	(g34917,I33143);
	not 	XG20647 	(g34919,I33149);
	not 	XG20648 	(g34921,I33155);
	not 	XG20649 	(g34923,I33161);
	not 	XG20650 	(g34925,I33167);
	not 	XG20651 	(g34927,I33173);
	not 	XG20652 	(g34956,I33214);
	not 	XG20653 	(g34972,I33232);
	not 	XG20654 	(g24168,I23348);
	not 	XG20655 	(g24178,I23378);
	not 	XG20656 	(g12833,I15448);
	not 	XG20657 	(g24174,I23366);
	not 	XG20658 	(g24181,I23387);
	not 	XG20659 	(g24172,I23360);
	not 	XG20660 	(g24161,I23327);
	not 	XG20661 	(g24177,I23375);
	not 	XG20662 	(g24171,I23357);
	not 	XG20663 	(g24163,I23333);
	not 	XG20664 	(g24170,I23354);
	not 	XG20665 	(g24185,I23399);
	not 	XG20666 	(g24164,I23336);
	not 	XG20667 	(g24173,I23363);
	not 	XG20668 	(g24162,I23330);
	not 	XG20669 	(g24179,I23381);
	not 	XG20670 	(g24180,I23384);
	not 	XG20671 	(g24175,I23369);
	not 	XG20672 	(g24183,I23393);
	not 	XG20673 	(g24166,I23342);
	not 	XG20674 	(g24176,I23372);
	not 	XG20675 	(g24184,I23396);
	not 	XG20676 	(g24169,I23351);
	not 	XG20677 	(g24182,I23390);
	not 	XG20678 	(g24165,I23339);
	not 	XG20679 	(g24167,I23345);

endmodule

